magic
tech sky130A
magscale 1 2
timestamp 1656242432
<< viali >>
rect 17049 20553 17083 20587
rect 14749 20485 14783 20519
rect 5825 20417 5859 20451
rect 6377 20417 6411 20451
rect 8401 20417 8435 20451
rect 9045 20417 9079 20451
rect 12642 20417 12676 20451
rect 15853 20417 15887 20451
rect 16129 20417 16163 20451
rect 17233 20417 17267 20451
rect 17509 20417 17543 20451
rect 18061 20417 18095 20451
rect 18613 20417 18647 20451
rect 20085 20417 20119 20451
rect 20545 20417 20579 20451
rect 8125 20349 8159 20383
rect 9505 20349 9539 20383
rect 12909 20349 12943 20383
rect 15485 20349 15519 20383
rect 19809 20349 19843 20383
rect 21189 20349 21223 20383
rect 8585 20281 8619 20315
rect 17693 20281 17727 20315
rect 6009 20213 6043 20247
rect 9229 20213 9263 20247
rect 11529 20213 11563 20247
rect 13277 20213 13311 20247
rect 15117 20213 15151 20247
rect 16313 20213 16347 20247
rect 18245 20213 18279 20247
rect 18797 20213 18831 20247
rect 8953 20009 8987 20043
rect 13093 20009 13127 20043
rect 16037 20009 16071 20043
rect 8585 19941 8619 19975
rect 15393 19941 15427 19975
rect 8033 19873 8067 19907
rect 9597 19873 9631 19907
rect 18797 19873 18831 19907
rect 21373 19873 21407 19907
rect 8217 19805 8251 19839
rect 10425 19805 10459 19839
rect 11345 19805 11379 19839
rect 13369 19805 13403 19839
rect 14749 19805 14783 19839
rect 15209 19805 15243 19839
rect 16313 19805 16347 19839
rect 16773 19805 16807 19839
rect 19441 19805 19475 19839
rect 9321 19737 9355 19771
rect 9965 19737 9999 19771
rect 11590 19737 11624 19771
rect 18552 19737 18586 19771
rect 21128 19737 21162 19771
rect 7573 19669 7607 19703
rect 8125 19669 8159 19703
rect 9413 19669 9447 19703
rect 10609 19669 10643 19703
rect 12725 19669 12759 19703
rect 13553 19669 13587 19703
rect 14933 19669 14967 19703
rect 16497 19669 16531 19703
rect 16957 19669 16991 19703
rect 17417 19669 17451 19703
rect 19625 19669 19659 19703
rect 19993 19669 20027 19703
rect 7113 19465 7147 19499
rect 7389 19465 7423 19499
rect 7757 19465 7791 19499
rect 8769 19465 8803 19499
rect 13645 19465 13679 19499
rect 18613 19465 18647 19499
rect 8861 19397 8895 19431
rect 10894 19397 10928 19431
rect 12510 19397 12544 19431
rect 15178 19397 15212 19431
rect 6929 19329 6963 19363
rect 7849 19329 7883 19363
rect 17489 19329 17523 19363
rect 19145 19329 19179 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 8033 19261 8067 19295
rect 9045 19261 9079 19295
rect 11161 19261 11195 19295
rect 11529 19261 11563 19295
rect 12265 19261 12299 19295
rect 14933 19261 14967 19295
rect 17233 19261 17267 19295
rect 18889 19261 18923 19295
rect 9781 19193 9815 19227
rect 8401 19125 8435 19159
rect 13921 19125 13955 19159
rect 14565 19125 14599 19159
rect 16313 19125 16347 19159
rect 16773 19125 16807 19159
rect 20269 19125 20303 19159
rect 20729 19125 20763 19159
rect 21281 19125 21315 19159
rect 11253 18921 11287 18955
rect 8217 18717 8251 18751
rect 9873 18717 9907 18751
rect 12909 18717 12943 18751
rect 14289 18717 14323 18751
rect 14556 18717 14590 18751
rect 17325 18717 17359 18751
rect 18705 18717 18739 18751
rect 19257 18717 19291 18751
rect 21097 18717 21131 18751
rect 10140 18649 10174 18683
rect 12642 18649 12676 18683
rect 17080 18649 17114 18683
rect 19524 18649 19558 18683
rect 8401 18581 8435 18615
rect 9321 18581 9355 18615
rect 11529 18581 11563 18615
rect 13277 18581 13311 18615
rect 15669 18581 15703 18615
rect 15945 18581 15979 18615
rect 17693 18581 17727 18615
rect 17969 18581 18003 18615
rect 18337 18581 18371 18615
rect 18889 18581 18923 18615
rect 20637 18581 20671 18615
rect 21281 18581 21315 18615
rect 8861 18377 8895 18411
rect 9229 18377 9263 18411
rect 11529 18377 11563 18411
rect 12081 18377 12115 18411
rect 18981 18377 19015 18411
rect 13194 18241 13228 18275
rect 16057 18241 16091 18275
rect 17132 18241 17166 18275
rect 19165 18241 19199 18275
rect 19441 18241 19475 18275
rect 20260 18241 20294 18275
rect 9321 18173 9355 18207
rect 9505 18173 9539 18207
rect 13461 18173 13495 18207
rect 16313 18173 16347 18207
rect 16865 18173 16899 18207
rect 19993 18173 20027 18207
rect 14933 18105 14967 18139
rect 18521 18105 18555 18139
rect 19625 18105 19659 18139
rect 13737 18037 13771 18071
rect 14565 18037 14599 18071
rect 18245 18037 18279 18071
rect 21373 18037 21407 18071
rect 18889 17833 18923 17867
rect 16497 17765 16531 17799
rect 12918 17629 12952 17663
rect 13185 17629 13219 17663
rect 17621 17629 17655 17663
rect 17877 17629 17911 17663
rect 18153 17629 18187 17663
rect 18705 17629 18739 17663
rect 20637 17629 20671 17663
rect 21097 17629 21131 17663
rect 20370 17561 20404 17595
rect 11805 17493 11839 17527
rect 13461 17493 13495 17527
rect 15025 17493 15059 17527
rect 15393 17493 15427 17527
rect 15761 17493 15795 17527
rect 16129 17493 16163 17527
rect 19257 17493 19291 17527
rect 21281 17493 21315 17527
rect 11713 17289 11747 17323
rect 16681 17221 16715 17255
rect 12081 17153 12115 17187
rect 12348 17153 12382 17187
rect 15200 17153 15234 17187
rect 18357 17153 18391 17187
rect 18613 17153 18647 17187
rect 19165 17153 19199 17187
rect 19708 17153 19742 17187
rect 21097 17153 21131 17187
rect 14933 17085 14967 17119
rect 19441 17085 19475 17119
rect 13737 17017 13771 17051
rect 16313 17017 16347 17051
rect 18981 17017 19015 17051
rect 21281 17017 21315 17051
rect 13461 16949 13495 16983
rect 17233 16949 17267 16983
rect 20821 16949 20855 16983
rect 10517 16745 10551 16779
rect 9965 16677 9999 16711
rect 9413 16609 9447 16643
rect 9597 16609 9631 16643
rect 11897 16609 11931 16643
rect 12173 16609 12207 16643
rect 14289 16609 14323 16643
rect 11641 16541 11675 16575
rect 15945 16541 15979 16575
rect 17601 16541 17635 16575
rect 17969 16541 18003 16575
rect 18337 16541 18371 16575
rect 18705 16541 18739 16575
rect 20637 16541 20671 16575
rect 21097 16541 21131 16575
rect 9321 16473 9355 16507
rect 12418 16473 12452 16507
rect 14556 16473 14590 16507
rect 16212 16473 16246 16507
rect 20392 16473 20426 16507
rect 8493 16405 8527 16439
rect 8953 16405 8987 16439
rect 13553 16405 13587 16439
rect 15669 16405 15703 16439
rect 17325 16405 17359 16439
rect 18889 16405 18923 16439
rect 19257 16405 19291 16439
rect 21281 16405 21315 16439
rect 15853 16201 15887 16235
rect 19441 16201 19475 16235
rect 12642 16065 12676 16099
rect 17805 16065 17839 16099
rect 19625 16065 19659 16099
rect 20157 16065 20191 16099
rect 12909 15997 12943 16031
rect 18061 15997 18095 16031
rect 18337 15997 18371 16031
rect 18981 15997 19015 16031
rect 19901 15997 19935 16031
rect 11529 15861 11563 15895
rect 13277 15861 13311 15895
rect 13645 15861 13679 15895
rect 16681 15861 16715 15895
rect 21281 15861 21315 15895
rect 15853 15521 15887 15555
rect 16129 15521 16163 15555
rect 16497 15521 16531 15555
rect 17049 15521 17083 15555
rect 17417 15521 17451 15555
rect 17785 15521 17819 15555
rect 18153 15521 18187 15555
rect 18797 15521 18831 15555
rect 12449 15453 12483 15487
rect 19717 15453 19751 15487
rect 21373 15453 21407 15487
rect 12182 15385 12216 15419
rect 15608 15385 15642 15419
rect 21128 15385 21162 15419
rect 11069 15317 11103 15351
rect 12817 15317 12851 15351
rect 14473 15317 14507 15351
rect 19533 15317 19567 15351
rect 19993 15317 20027 15351
rect 16313 15113 16347 15147
rect 17805 15045 17839 15079
rect 13021 14977 13055 15011
rect 14832 14977 14866 15011
rect 18061 14977 18095 15011
rect 19461 14977 19495 15011
rect 19717 14977 19751 15011
rect 21117 14977 21151 15011
rect 21373 14977 21407 15011
rect 13277 14909 13311 14943
rect 14565 14909 14599 14943
rect 15945 14841 15979 14875
rect 11897 14773 11931 14807
rect 13645 14773 13679 14807
rect 16681 14773 16715 14807
rect 18337 14773 18371 14807
rect 19993 14773 20027 14807
rect 19533 14569 19567 14603
rect 16129 14501 16163 14535
rect 12081 14365 12115 14399
rect 13737 14365 13771 14399
rect 14105 14365 14139 14399
rect 14473 14365 14507 14399
rect 17509 14365 17543 14399
rect 17785 14365 17819 14399
rect 18337 14365 18371 14399
rect 18797 14365 18831 14399
rect 19717 14365 19751 14399
rect 21373 14365 21407 14399
rect 11836 14297 11870 14331
rect 13492 14297 13526 14331
rect 14740 14297 14774 14331
rect 17253 14297 17287 14331
rect 21106 14297 21140 14331
rect 10701 14229 10735 14263
rect 12357 14229 12391 14263
rect 15853 14229 15887 14263
rect 19993 14229 20027 14263
rect 8677 14025 8711 14059
rect 13369 14025 13403 14059
rect 18245 14025 18279 14059
rect 19901 14025 19935 14059
rect 20729 14025 20763 14059
rect 8217 13957 8251 13991
rect 9045 13957 9079 13991
rect 17132 13957 17166 13991
rect 18788 13957 18822 13991
rect 8309 13889 8343 13923
rect 12256 13889 12290 13923
rect 16865 13889 16899 13923
rect 18521 13889 18555 13923
rect 20545 13889 20579 13923
rect 21097 13889 21131 13923
rect 8125 13821 8159 13855
rect 11989 13821 12023 13855
rect 16037 13821 16071 13855
rect 11621 13685 11655 13719
rect 13645 13685 13679 13719
rect 20177 13685 20211 13719
rect 21281 13685 21315 13719
rect 21373 13481 21407 13515
rect 11161 13345 11195 13379
rect 15669 13345 15703 13379
rect 18429 13345 18463 13379
rect 18705 13345 18739 13379
rect 19993 13345 20027 13379
rect 12817 13277 12851 13311
rect 15945 13277 15979 13311
rect 19533 13277 19567 13311
rect 20249 13277 20283 13311
rect 11428 13209 11462 13243
rect 18162 13209 18196 13243
rect 12541 13141 12575 13175
rect 15853 13141 15887 13175
rect 16313 13141 16347 13175
rect 16589 13141 16623 13175
rect 17049 13141 17083 13175
rect 19717 13141 19751 13175
rect 15485 12937 15519 12971
rect 18705 12937 18739 12971
rect 20821 12937 20855 12971
rect 21281 12937 21315 12971
rect 17509 12869 17543 12903
rect 15117 12801 15151 12835
rect 15761 12801 15795 12835
rect 17417 12801 17451 12835
rect 18061 12801 18095 12835
rect 19073 12801 19107 12835
rect 19717 12801 19751 12835
rect 20177 12801 20211 12835
rect 20637 12801 20671 12835
rect 21097 12801 21131 12835
rect 14841 12733 14875 12767
rect 15025 12733 15059 12767
rect 17601 12733 17635 12767
rect 19165 12733 19199 12767
rect 19349 12733 19383 12767
rect 17049 12665 17083 12699
rect 12909 12597 12943 12631
rect 16773 12597 16807 12631
rect 20361 12597 20395 12631
rect 11989 12393 12023 12427
rect 14841 12393 14875 12427
rect 16313 12393 16347 12427
rect 19257 12393 19291 12427
rect 20637 12393 20671 12427
rect 21281 12393 21315 12427
rect 10517 12325 10551 12359
rect 18797 12325 18831 12359
rect 9873 12257 9907 12291
rect 10057 12257 10091 12291
rect 12541 12257 12575 12291
rect 13553 12257 13587 12291
rect 14197 12257 14231 12291
rect 15853 12257 15887 12291
rect 16865 12257 16899 12291
rect 17877 12257 17911 12291
rect 19901 12257 19935 12291
rect 12449 12189 12483 12223
rect 14381 12189 14415 12223
rect 15669 12189 15703 12223
rect 16773 12189 16807 12223
rect 18337 12189 18371 12223
rect 19625 12189 19659 12223
rect 20821 12189 20855 12223
rect 21097 12189 21131 12223
rect 10149 12121 10183 12155
rect 10793 12121 10827 12155
rect 14473 12121 14507 12155
rect 15761 12121 15795 12155
rect 20269 12121 20303 12155
rect 11621 12053 11655 12087
rect 12357 12053 12391 12087
rect 13001 12053 13035 12087
rect 13369 12053 13403 12087
rect 13461 12053 13495 12087
rect 15301 12053 15335 12087
rect 16681 12053 16715 12087
rect 17325 12053 17359 12087
rect 17693 12053 17727 12087
rect 17785 12053 17819 12087
rect 18521 12053 18555 12087
rect 19717 12053 19751 12087
rect 11989 11849 12023 11883
rect 15301 11849 15335 11883
rect 17693 11849 17727 11883
rect 18245 11849 18279 11883
rect 19257 11849 19291 11883
rect 19717 11849 19751 11883
rect 20453 11849 20487 11883
rect 21189 11849 21223 11883
rect 2053 11781 2087 11815
rect 1685 11713 1719 11747
rect 11713 11713 11747 11747
rect 12357 11713 12391 11747
rect 14933 11713 14967 11747
rect 15577 11713 15611 11747
rect 16681 11713 16715 11747
rect 17601 11713 17635 11747
rect 18613 11713 18647 11747
rect 19625 11713 19659 11747
rect 20269 11713 20303 11747
rect 20913 11713 20947 11747
rect 21373 11713 21407 11747
rect 12449 11645 12483 11679
rect 12633 11645 12667 11679
rect 14657 11645 14691 11679
rect 14841 11645 14875 11679
rect 17785 11645 17819 11679
rect 18705 11645 18739 11679
rect 18797 11645 18831 11679
rect 19901 11645 19935 11679
rect 20729 11577 20763 11611
rect 1501 11509 1535 11543
rect 16129 11509 16163 11543
rect 16865 11509 16899 11543
rect 17233 11509 17267 11543
rect 14933 11305 14967 11339
rect 17325 11305 17359 11339
rect 17785 11305 17819 11339
rect 18705 11305 18739 11339
rect 19533 11305 19567 11339
rect 19809 11305 19843 11339
rect 20269 11305 20303 11339
rect 20729 11305 20763 11339
rect 21189 11305 21223 11339
rect 14289 11169 14323 11203
rect 14473 11169 14507 11203
rect 16037 11169 16071 11203
rect 18061 11169 18095 11203
rect 17141 11101 17175 11135
rect 17601 11101 17635 11135
rect 18889 11101 18923 11135
rect 19349 11101 19383 11135
rect 19993 11101 20027 11135
rect 20453 11101 20487 11135
rect 20913 11101 20947 11135
rect 21373 11101 21407 11135
rect 14565 11033 14599 11067
rect 16405 11033 16439 11067
rect 15301 10965 15335 10999
rect 16681 10965 16715 10999
rect 15209 10761 15243 10795
rect 15577 10761 15611 10795
rect 17693 10761 17727 10795
rect 18153 10761 18187 10795
rect 18613 10761 18647 10795
rect 20085 10761 20119 10795
rect 20545 10761 20579 10795
rect 21005 10761 21039 10795
rect 21373 10761 21407 10795
rect 17325 10625 17359 10659
rect 17969 10625 18003 10659
rect 18429 10625 18463 10659
rect 18889 10625 18923 10659
rect 19441 10625 19475 10659
rect 19901 10625 19935 10659
rect 20361 10625 20395 10659
rect 20821 10625 20855 10659
rect 14933 10557 14967 10591
rect 15117 10557 15151 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 19073 10489 19107 10523
rect 19625 10421 19659 10455
rect 15025 10217 15059 10251
rect 17049 10217 17083 10251
rect 18705 10217 18739 10251
rect 19625 10217 19659 10251
rect 20085 10149 20119 10183
rect 20361 10149 20395 10183
rect 15577 10081 15611 10115
rect 16497 10081 16531 10115
rect 18061 10081 18095 10115
rect 21005 10081 21039 10115
rect 15485 10013 15519 10047
rect 16681 10013 16715 10047
rect 17693 10013 17727 10047
rect 19441 10013 19475 10047
rect 19901 10013 19935 10047
rect 15393 9945 15427 9979
rect 16589 9945 16623 9979
rect 14749 9877 14783 9911
rect 17509 9877 17543 9911
rect 18245 9877 18279 9911
rect 18337 9877 18371 9911
rect 20729 9877 20763 9911
rect 20821 9877 20855 9911
rect 17509 9673 17543 9707
rect 18245 9673 18279 9707
rect 18705 9673 18739 9707
rect 19717 9673 19751 9707
rect 20177 9673 20211 9707
rect 15209 9605 15243 9639
rect 12541 9537 12575 9571
rect 17785 9537 17819 9571
rect 18613 9537 18647 9571
rect 19533 9537 19567 9571
rect 20545 9537 20579 9571
rect 21373 9537 21407 9571
rect 12633 9469 12667 9503
rect 12725 9469 12759 9503
rect 14933 9469 14967 9503
rect 15117 9469 15151 9503
rect 18797 9469 18831 9503
rect 20637 9469 20671 9503
rect 20821 9469 20855 9503
rect 12173 9401 12207 9435
rect 17969 9401 18003 9435
rect 15577 9333 15611 9367
rect 17141 9333 17175 9367
rect 21189 9333 21223 9367
rect 15577 9129 15611 9163
rect 16957 9129 16991 9163
rect 17969 9129 18003 9163
rect 19349 9129 19383 9163
rect 20821 9129 20855 9163
rect 21097 9129 21131 9163
rect 19809 9061 19843 9095
rect 15025 8993 15059 9027
rect 16313 8993 16347 9027
rect 17417 8993 17451 9027
rect 20177 8993 20211 9027
rect 15853 8925 15887 8959
rect 16497 8925 16531 8959
rect 18889 8925 18923 8959
rect 19625 8925 19659 8959
rect 21281 8925 21315 8959
rect 15209 8857 15243 8891
rect 17601 8857 17635 8891
rect 18245 8857 18279 8891
rect 15117 8789 15151 8823
rect 16589 8789 16623 8823
rect 17509 8789 17543 8823
rect 18705 8789 18739 8823
rect 20361 8789 20395 8823
rect 20453 8789 20487 8823
rect 16313 8585 16347 8619
rect 17969 8585 18003 8619
rect 18429 8585 18463 8619
rect 19717 8585 19751 8619
rect 20729 8585 20763 8619
rect 21189 8585 21223 8619
rect 20085 8517 20119 8551
rect 16681 8449 16715 8483
rect 17233 8449 17267 8483
rect 17693 8449 17727 8483
rect 18337 8449 18371 8483
rect 19441 8449 19475 8483
rect 21373 8449 21407 8483
rect 18521 8381 18555 8415
rect 20177 8381 20211 8415
rect 20361 8381 20395 8415
rect 17509 8313 17543 8347
rect 19257 8313 19291 8347
rect 17693 8041 17727 8075
rect 20361 8041 20395 8075
rect 17049 7973 17083 8007
rect 18245 7905 18279 7939
rect 19533 7905 19567 7939
rect 21005 7905 21039 7939
rect 17417 7837 17451 7871
rect 18889 7837 18923 7871
rect 20821 7837 20855 7871
rect 18061 7769 18095 7803
rect 19625 7769 19659 7803
rect 20729 7769 20763 7803
rect 18153 7701 18187 7735
rect 18705 7701 18739 7735
rect 19717 7701 19751 7735
rect 20085 7701 20119 7735
rect 17049 7497 17083 7531
rect 19349 7497 19383 7531
rect 20361 7497 20395 7531
rect 20729 7497 20763 7531
rect 19625 7429 19659 7463
rect 17877 7361 17911 7395
rect 18337 7361 18371 7395
rect 18981 7361 19015 7395
rect 20269 7361 20303 7395
rect 21373 7361 21407 7395
rect 18705 7293 18739 7327
rect 18889 7293 18923 7327
rect 20177 7293 20211 7327
rect 16773 7225 16807 7259
rect 17509 7157 17543 7191
rect 18153 7157 18187 7191
rect 21189 7157 21223 7191
rect 16865 6817 16899 6851
rect 18061 6817 18095 6851
rect 18245 6817 18279 6851
rect 19901 6817 19935 6851
rect 20729 6817 20763 6851
rect 20913 6817 20947 6851
rect 17141 6749 17175 6783
rect 18705 6749 18739 6783
rect 19717 6749 19751 6783
rect 17969 6681 18003 6715
rect 19625 6681 19659 6715
rect 21373 6681 21407 6715
rect 17325 6613 17359 6647
rect 17601 6613 17635 6647
rect 18889 6613 18923 6647
rect 19257 6613 19291 6647
rect 20269 6613 20303 6647
rect 20637 6613 20671 6647
rect 18153 6409 18187 6443
rect 18521 6409 18555 6443
rect 20361 6409 20395 6443
rect 19625 6341 19659 6375
rect 20729 6341 20763 6375
rect 16957 6273 16991 6307
rect 17417 6273 17451 6307
rect 17877 6273 17911 6307
rect 20085 6273 20119 6307
rect 16313 6205 16347 6239
rect 18613 6205 18647 6239
rect 18705 6205 18739 6239
rect 20821 6205 20855 6239
rect 20913 6205 20947 6239
rect 17693 6137 17727 6171
rect 17233 6069 17267 6103
rect 19901 6069 19935 6103
rect 17601 5865 17635 5899
rect 19257 5865 19291 5899
rect 20453 5865 20487 5899
rect 17141 5797 17175 5831
rect 15669 5729 15703 5763
rect 19901 5729 19935 5763
rect 21005 5729 21039 5763
rect 16405 5661 16439 5695
rect 16865 5661 16899 5695
rect 17325 5661 17359 5695
rect 17785 5661 17819 5695
rect 18429 5661 18463 5695
rect 20821 5661 20855 5695
rect 16037 5593 16071 5627
rect 19625 5593 19659 5627
rect 16681 5525 16715 5559
rect 18245 5525 18279 5559
rect 18889 5525 18923 5559
rect 19717 5525 19751 5559
rect 20913 5525 20947 5559
rect 15853 5321 15887 5355
rect 16313 5321 16347 5355
rect 17141 5321 17175 5355
rect 19809 5321 19843 5355
rect 20177 5321 20211 5355
rect 15301 5253 15335 5287
rect 20821 5253 20855 5287
rect 15945 5185 15979 5219
rect 17049 5185 17083 5219
rect 17693 5185 17727 5219
rect 18981 5185 19015 5219
rect 19717 5185 19751 5219
rect 15761 5117 15795 5151
rect 17325 5117 17359 5151
rect 18337 5117 18371 5151
rect 19625 5117 19659 5151
rect 20913 5117 20947 5151
rect 21097 5117 21131 5151
rect 20453 5049 20487 5083
rect 16681 4981 16715 5015
rect 18797 4981 18831 5015
rect 16957 4777 16991 4811
rect 21281 4777 21315 4811
rect 16497 4709 16531 4743
rect 19993 4709 20027 4743
rect 14289 4641 14323 4675
rect 15945 4641 15979 4675
rect 18337 4641 18371 4675
rect 19441 4641 19475 4675
rect 20821 4641 20855 4675
rect 7297 4573 7331 4607
rect 14657 4573 14691 4607
rect 15485 4573 15519 4607
rect 16681 4573 16715 4607
rect 17141 4573 17175 4607
rect 17601 4573 17635 4607
rect 15209 4505 15243 4539
rect 18521 4505 18555 4539
rect 19625 4505 19659 4539
rect 20729 4505 20763 4539
rect 7481 4437 7515 4471
rect 15669 4437 15703 4471
rect 17417 4437 17451 4471
rect 18429 4437 18463 4471
rect 18889 4437 18923 4471
rect 19533 4437 19567 4471
rect 20269 4437 20303 4471
rect 20637 4437 20671 4471
rect 18245 4233 18279 4267
rect 19349 4233 19383 4267
rect 19441 4233 19475 4267
rect 14289 4097 14323 4131
rect 14749 4097 14783 4131
rect 15393 4097 15427 4131
rect 15669 4097 15703 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 17141 4097 17175 4131
rect 19993 4097 20027 4131
rect 14013 4029 14047 4063
rect 17969 4029 18003 4063
rect 18153 4029 18187 4063
rect 19533 4029 19567 4063
rect 20545 4029 20579 4063
rect 20821 4029 20855 4063
rect 18613 3961 18647 3995
rect 18981 3961 19015 3995
rect 20177 3961 20211 3995
rect 14473 3893 14507 3927
rect 14933 3893 14967 3927
rect 15209 3893 15243 3927
rect 15853 3893 15887 3927
rect 16313 3893 16347 3927
rect 16681 3893 16715 3927
rect 17325 3893 17359 3927
rect 16313 3689 16347 3723
rect 17601 3689 17635 3723
rect 18705 3689 18739 3723
rect 20269 3689 20303 3723
rect 14841 3621 14875 3655
rect 15485 3621 15519 3655
rect 17233 3621 17267 3655
rect 18061 3553 18095 3587
rect 18245 3553 18279 3587
rect 19717 3553 19751 3587
rect 19809 3553 19843 3587
rect 20821 3553 20855 3587
rect 13553 3485 13587 3519
rect 14381 3485 14415 3519
rect 15025 3485 15059 3519
rect 15301 3485 15335 3519
rect 16129 3485 16163 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 20545 3485 20579 3519
rect 13277 3417 13311 3451
rect 15853 3417 15887 3451
rect 18797 3417 18831 3451
rect 19901 3417 19935 3451
rect 3065 3349 3099 3383
rect 4353 3349 4387 3383
rect 13737 3349 13771 3383
rect 14565 3349 14599 3383
rect 16589 3349 16623 3383
rect 17969 3349 18003 3383
rect 2789 3145 2823 3179
rect 9229 3145 9263 3179
rect 12541 3145 12575 3179
rect 2605 3009 2639 3043
rect 3985 3009 4019 3043
rect 9045 3009 9079 3043
rect 13185 3009 13219 3043
rect 13645 3009 13679 3043
rect 14105 3009 14139 3043
rect 14565 3009 14599 3043
rect 15209 3009 15243 3043
rect 15485 3009 15519 3043
rect 16221 3009 16255 3043
rect 17141 3009 17175 3043
rect 17693 3009 17727 3043
rect 18245 3009 18279 3043
rect 18797 3009 18831 3043
rect 19349 3009 19383 3043
rect 19901 3009 19935 3043
rect 20821 3009 20855 3043
rect 12909 2941 12943 2975
rect 20545 2941 20579 2975
rect 4169 2873 4203 2907
rect 14289 2873 14323 2907
rect 14749 2873 14783 2907
rect 17877 2873 17911 2907
rect 2329 2805 2363 2839
rect 3341 2805 3375 2839
rect 3709 2805 3743 2839
rect 4813 2805 4847 2839
rect 5273 2805 5307 2839
rect 5733 2805 5767 2839
rect 6377 2805 6411 2839
rect 6929 2805 6963 2839
rect 7205 2805 7239 2839
rect 7573 2805 7607 2839
rect 8033 2805 8067 2839
rect 8401 2805 8435 2839
rect 8677 2805 8711 2839
rect 9505 2805 9539 2839
rect 9873 2805 9907 2839
rect 10333 2805 10367 2839
rect 10793 2805 10827 2839
rect 11529 2805 11563 2839
rect 13369 2805 13403 2839
rect 13829 2805 13863 2839
rect 15025 2805 15059 2839
rect 15669 2805 15703 2839
rect 16037 2805 16071 2839
rect 16957 2805 16991 2839
rect 18429 2805 18463 2839
rect 18981 2805 19015 2839
rect 19533 2805 19567 2839
rect 20085 2805 20119 2839
rect 5089 2601 5123 2635
rect 7205 2601 7239 2635
rect 7665 2601 7699 2635
rect 8125 2601 8159 2635
rect 8585 2601 8619 2635
rect 9781 2601 9815 2635
rect 11161 2601 11195 2635
rect 15945 2601 15979 2635
rect 4169 2533 4203 2567
rect 6009 2533 6043 2567
rect 9321 2533 9355 2567
rect 14749 2533 14783 2567
rect 17969 2533 18003 2567
rect 19993 2465 20027 2499
rect 20821 2465 20855 2499
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 3985 2397 4019 2431
rect 4445 2397 4479 2431
rect 4905 2397 4939 2431
rect 5365 2397 5399 2431
rect 5825 2397 5859 2431
rect 6561 2397 6595 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 9597 2397 9631 2431
rect 10057 2397 10091 2431
rect 10517 2397 10551 2431
rect 10977 2397 11011 2431
rect 11897 2397 11931 2431
rect 12449 2397 12483 2431
rect 13001 2397 13035 2431
rect 13553 2397 13587 2431
rect 14381 2397 14415 2431
rect 14933 2397 14967 2431
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 17785 2397 17819 2431
rect 18613 2397 18647 2431
rect 20269 2397 20303 2431
rect 20545 2397 20579 2431
rect 2237 2329 2271 2363
rect 1869 2261 1903 2295
rect 2329 2261 2363 2295
rect 2973 2261 3007 2295
rect 3433 2261 3467 2295
rect 4629 2261 4663 2295
rect 5549 2261 5583 2295
rect 6745 2261 6779 2295
rect 10241 2261 10275 2295
rect 10701 2261 10735 2295
rect 11713 2261 11747 2295
rect 12265 2261 12299 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 14197 2261 14231 2295
rect 15301 2261 15335 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 18429 2261 18463 2295
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 18046 20584 18052 20596
rect 17083 20556 18052 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 19306 20556 20576 20584
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 14737 20519 14795 20525
rect 7156 20488 14412 20516
rect 7156 20476 7162 20488
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5776 20420 5825 20448
rect 5776 20408 5782 20420
rect 5813 20417 5825 20420
rect 5859 20448 5871 20451
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 5859 20420 6377 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 8389 20451 8447 20457
rect 8389 20417 8401 20451
rect 8435 20448 8447 20451
rect 8570 20448 8576 20460
rect 8435 20420 8576 20448
rect 8435 20417 8447 20420
rect 8389 20411 8447 20417
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 9033 20451 9091 20457
rect 9033 20417 9045 20451
rect 9079 20448 9091 20451
rect 9122 20448 9128 20460
rect 9079 20420 9128 20448
rect 9079 20417 9091 20420
rect 9033 20411 9091 20417
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 12630 20451 12688 20457
rect 12630 20448 12642 20451
rect 11756 20420 12642 20448
rect 11756 20408 11762 20420
rect 12630 20417 12642 20420
rect 12676 20417 12688 20451
rect 14384 20448 14412 20488
rect 14737 20485 14749 20519
rect 14783 20516 14795 20519
rect 19306 20516 19334 20556
rect 14783 20488 19334 20516
rect 14783 20485 14795 20488
rect 14737 20479 14795 20485
rect 15286 20448 15292 20460
rect 14384 20420 15292 20448
rect 12630 20411 12688 20417
rect 15286 20408 15292 20420
rect 15344 20408 15350 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 15887 20420 16129 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16117 20417 16129 20420
rect 16163 20448 16175 20451
rect 17126 20448 17132 20460
rect 16163 20420 17132 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20448 17279 20451
rect 17310 20448 17316 20460
rect 17267 20420 17316 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 17310 20408 17316 20420
rect 17368 20408 17374 20460
rect 17494 20448 17500 20460
rect 17455 20420 17500 20448
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17644 20420 18061 20448
rect 17644 20408 17650 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 18196 20420 18613 20448
rect 18196 20408 18202 20420
rect 18601 20417 18613 20420
rect 18647 20417 18659 20451
rect 20070 20448 20076 20460
rect 18601 20411 18659 20417
rect 19260 20420 20076 20448
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 8202 20380 8208 20392
rect 8159 20352 8208 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 9490 20380 9496 20392
rect 9451 20352 9496 20380
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20380 12955 20383
rect 15473 20383 15531 20389
rect 12943 20352 13308 20380
rect 12943 20349 12955 20352
rect 12897 20343 12955 20349
rect 8573 20315 8631 20321
rect 8573 20281 8585 20315
rect 8619 20312 8631 20315
rect 13170 20312 13176 20324
rect 8619 20284 12020 20312
rect 8619 20281 8631 20284
rect 8573 20275 8631 20281
rect 5994 20244 6000 20256
rect 5955 20216 6000 20244
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 9214 20244 9220 20256
rect 9175 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9582 20204 9588 20256
rect 9640 20244 9646 20256
rect 10870 20244 10876 20256
rect 9640 20216 10876 20244
rect 9640 20204 9646 20216
rect 10870 20204 10876 20216
rect 10928 20244 10934 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 10928 20216 11529 20244
rect 10928 20204 10934 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11992 20244 12020 20284
rect 13004 20284 13176 20312
rect 13004 20244 13032 20284
rect 13170 20272 13176 20284
rect 13228 20272 13234 20324
rect 11992 20216 13032 20244
rect 11517 20207 11575 20213
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13280 20253 13308 20352
rect 15473 20349 15485 20383
rect 15519 20380 15531 20383
rect 19260 20380 19288 20420
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20548 20457 20576 20556
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20622 20448 20628 20460
rect 20579 20420 20628 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 15519 20352 19288 20380
rect 19797 20383 19855 20389
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 19797 20349 19809 20383
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21358 20380 21364 20392
rect 21223 20352 21364 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 17681 20315 17739 20321
rect 17681 20281 17693 20315
rect 17727 20312 17739 20315
rect 17954 20312 17960 20324
rect 17727 20284 17960 20312
rect 17727 20281 17739 20284
rect 17681 20275 17739 20281
rect 17954 20272 17960 20284
rect 18012 20272 18018 20324
rect 19812 20312 19840 20343
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 22462 20312 22468 20324
rect 19812 20284 22468 20312
rect 22462 20272 22468 20284
rect 22520 20272 22526 20324
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 13136 20216 13277 20244
rect 13136 20204 13142 20216
rect 13265 20213 13277 20216
rect 13311 20244 13323 20247
rect 15102 20244 15108 20256
rect 13311 20216 15108 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 16301 20247 16359 20253
rect 16301 20213 16313 20247
rect 16347 20244 16359 20247
rect 18046 20244 18052 20256
rect 16347 20216 18052 20244
rect 16347 20213 16359 20216
rect 16301 20207 16359 20213
rect 18046 20204 18052 20216
rect 18104 20204 18110 20256
rect 18230 20244 18236 20256
rect 18191 20216 18236 20244
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 18782 20244 18788 20256
rect 18743 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 8941 20043 8999 20049
rect 8941 20009 8953 20043
rect 8987 20040 8999 20043
rect 9122 20040 9128 20052
rect 8987 20012 9128 20040
rect 8987 20009 8999 20012
rect 8941 20003 8999 20009
rect 9122 20000 9128 20012
rect 9180 20000 9186 20052
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 13078 20040 13084 20052
rect 9272 20012 12434 20040
rect 13039 20012 13084 20040
rect 9272 20000 9278 20012
rect 8573 19975 8631 19981
rect 8573 19941 8585 19975
rect 8619 19972 8631 19975
rect 12406 19972 12434 20012
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 15102 20000 15108 20052
rect 15160 20040 15166 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15160 20012 16037 20040
rect 15160 20000 15166 20012
rect 16025 20009 16037 20012
rect 16071 20040 16083 20043
rect 16071 20012 18828 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 15381 19975 15439 19981
rect 8619 19944 10456 19972
rect 12406 19944 15240 19972
rect 8619 19941 8631 19944
rect 8573 19935 8631 19941
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19904 8079 19907
rect 9398 19904 9404 19916
rect 8067 19876 9404 19904
rect 8067 19873 8079 19876
rect 8021 19867 8079 19873
rect 9398 19864 9404 19876
rect 9456 19864 9462 19916
rect 9582 19904 9588 19916
rect 9543 19876 9588 19904
rect 9582 19864 9588 19876
rect 9640 19864 9646 19916
rect 8202 19836 8208 19848
rect 8163 19808 8208 19836
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 10428 19845 10456 19944
rect 13170 19864 13176 19916
rect 13228 19904 13234 19916
rect 13228 19876 14780 19904
rect 13228 19864 13234 19876
rect 10413 19839 10471 19845
rect 10413 19805 10425 19839
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 11146 19796 11152 19848
rect 11204 19836 11210 19848
rect 11333 19839 11391 19845
rect 11333 19836 11345 19839
rect 11204 19808 11345 19836
rect 11204 19796 11210 19808
rect 11333 19805 11345 19808
rect 11379 19836 11391 19839
rect 13078 19836 13084 19848
rect 11379 19808 13084 19836
rect 11379 19805 11391 19808
rect 11333 19799 11391 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 14752 19845 14780 19876
rect 15212 19845 15240 19944
rect 15381 19941 15393 19975
rect 15427 19972 15439 19975
rect 17586 19972 17592 19984
rect 15427 19944 17592 19972
rect 15427 19941 15439 19944
rect 15381 19935 15439 19941
rect 17586 19932 17592 19944
rect 17644 19932 17650 19984
rect 17494 19904 17500 19916
rect 16408 19876 17500 19904
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 9953 19771 10011 19777
rect 9953 19768 9965 19771
rect 9355 19740 9965 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 9953 19737 9965 19740
rect 9999 19737 10011 19771
rect 9953 19731 10011 19737
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 11578 19771 11636 19777
rect 11578 19768 11590 19771
rect 11296 19740 11590 19768
rect 11296 19728 11302 19740
rect 11578 19737 11590 19740
rect 11624 19737 11636 19771
rect 13372 19768 13400 19799
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 16301 19839 16359 19845
rect 16301 19836 16313 19839
rect 15344 19808 16313 19836
rect 15344 19796 15350 19808
rect 16301 19805 16313 19808
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16408 19768 16436 19876
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 18800 19913 18828 20012
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 21358 19904 21364 19916
rect 18831 19876 19564 19904
rect 21319 19876 21364 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 16761 19839 16819 19845
rect 16761 19805 16773 19839
rect 16807 19836 16819 19839
rect 16850 19836 16856 19848
rect 16807 19808 16856 19836
rect 16807 19805 16819 19808
rect 16761 19799 16819 19805
rect 16850 19796 16856 19808
rect 16908 19796 16914 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 16960 19808 19441 19836
rect 11578 19731 11636 19737
rect 12406 19740 13400 19768
rect 13556 19740 16436 19768
rect 7561 19703 7619 19709
rect 7561 19669 7573 19703
rect 7607 19700 7619 19703
rect 7742 19700 7748 19712
rect 7607 19672 7748 19700
rect 7607 19669 7619 19672
rect 7561 19663 7619 19669
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 8113 19703 8171 19709
rect 8113 19669 8125 19703
rect 8159 19700 8171 19703
rect 8662 19700 8668 19712
rect 8159 19672 8668 19700
rect 8159 19669 8171 19672
rect 8113 19663 8171 19669
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19700 9459 19703
rect 10502 19700 10508 19712
rect 9447 19672 10508 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 10597 19703 10655 19709
rect 10597 19669 10609 19703
rect 10643 19700 10655 19703
rect 12406 19700 12434 19740
rect 10643 19672 12434 19700
rect 10643 19669 10655 19672
rect 10597 19663 10655 19669
rect 12618 19660 12624 19712
rect 12676 19700 12682 19712
rect 13556 19709 13584 19740
rect 12713 19703 12771 19709
rect 12713 19700 12725 19703
rect 12676 19672 12725 19700
rect 12676 19660 12682 19672
rect 12713 19669 12725 19672
rect 12759 19669 12771 19703
rect 12713 19663 12771 19669
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19669 13599 19703
rect 14918 19700 14924 19712
rect 14879 19672 14924 19700
rect 13541 19663 13599 19669
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 16390 19660 16396 19712
rect 16448 19700 16454 19712
rect 16960 19709 16988 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19536 19836 19564 19876
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 21376 19836 21404 19864
rect 19536 19808 21404 19836
rect 19429 19799 19487 19805
rect 18540 19771 18598 19777
rect 18540 19737 18552 19771
rect 18586 19768 18598 19771
rect 19702 19768 19708 19780
rect 18586 19740 19708 19768
rect 18586 19737 18598 19740
rect 18540 19731 18598 19737
rect 19702 19728 19708 19740
rect 19760 19728 19766 19780
rect 21116 19771 21174 19777
rect 21116 19737 21128 19771
rect 21162 19768 21174 19771
rect 21542 19768 21548 19780
rect 21162 19740 21548 19768
rect 21162 19737 21174 19740
rect 21116 19731 21174 19737
rect 21542 19728 21548 19740
rect 21600 19728 21606 19780
rect 16485 19703 16543 19709
rect 16485 19700 16497 19703
rect 16448 19672 16497 19700
rect 16448 19660 16454 19672
rect 16485 19669 16497 19672
rect 16531 19669 16543 19703
rect 16485 19663 16543 19669
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19669 17003 19703
rect 16945 19663 17003 19669
rect 17405 19703 17463 19709
rect 17405 19669 17417 19703
rect 17451 19700 17463 19703
rect 17586 19700 17592 19712
rect 17451 19672 17592 19700
rect 17451 19669 17463 19672
rect 17405 19663 17463 19669
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 19610 19700 19616 19712
rect 19571 19672 19616 19700
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 19981 19703 20039 19709
rect 19981 19669 19993 19703
rect 20027 19700 20039 19703
rect 20806 19700 20812 19712
rect 20027 19672 20812 19700
rect 20027 19669 20039 19672
rect 19981 19663 20039 19669
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 7098 19496 7104 19508
rect 7059 19468 7104 19496
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19465 7435 19499
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 7377 19459 7435 19465
rect 6917 19363 6975 19369
rect 6917 19329 6929 19363
rect 6963 19360 6975 19363
rect 7392 19360 7420 19459
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 9490 19496 9496 19508
rect 8803 19468 9496 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 10502 19456 10508 19508
rect 10560 19496 10566 19508
rect 11974 19496 11980 19508
rect 10560 19468 11980 19496
rect 10560 19456 10566 19468
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 13633 19499 13691 19505
rect 13633 19465 13645 19499
rect 13679 19465 13691 19499
rect 13633 19459 13691 19465
rect 8846 19428 8852 19440
rect 8807 19400 8852 19428
rect 8846 19388 8852 19400
rect 8904 19388 8910 19440
rect 9858 19388 9864 19440
rect 9916 19428 9922 19440
rect 10778 19428 10784 19440
rect 9916 19400 10784 19428
rect 9916 19388 9922 19400
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 10870 19388 10876 19440
rect 10928 19437 10934 19440
rect 10928 19428 10940 19437
rect 10928 19400 10973 19428
rect 10928 19391 10940 19400
rect 10928 19388 10934 19391
rect 11054 19388 11060 19440
rect 11112 19428 11118 19440
rect 12498 19431 12556 19437
rect 12498 19428 12510 19431
rect 11112 19400 12510 19428
rect 11112 19388 11118 19400
rect 12498 19397 12510 19400
rect 12544 19397 12556 19431
rect 12498 19391 12556 19397
rect 13648 19428 13676 19459
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 18138 19496 18144 19508
rect 14976 19468 18144 19496
rect 14976 19456 14982 19468
rect 18138 19456 18144 19468
rect 18196 19456 18202 19508
rect 18506 19456 18512 19508
rect 18564 19496 18570 19508
rect 18601 19499 18659 19505
rect 18601 19496 18613 19499
rect 18564 19468 18613 19496
rect 18564 19456 18570 19468
rect 18601 19465 18613 19468
rect 18647 19465 18659 19499
rect 18601 19459 18659 19465
rect 18874 19456 18880 19508
rect 18932 19496 18938 19508
rect 18932 19468 21128 19496
rect 18932 19456 18938 19468
rect 15166 19431 15224 19437
rect 15166 19428 15178 19431
rect 13648 19400 15178 19428
rect 6963 19332 7420 19360
rect 6963 19329 6975 19332
rect 6917 19323 6975 19329
rect 7834 19320 7840 19372
rect 7892 19360 7898 19372
rect 7892 19332 7937 19360
rect 7892 19320 7898 19332
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 13648 19360 13676 19400
rect 15166 19397 15178 19400
rect 15212 19397 15224 19431
rect 15166 19391 15224 19397
rect 16390 19388 16396 19440
rect 16448 19428 16454 19440
rect 16448 19400 20576 19428
rect 16448 19388 16454 19400
rect 17477 19363 17535 19369
rect 17477 19360 17489 19363
rect 9456 19332 13676 19360
rect 16592 19332 17489 19360
rect 9456 19320 9462 19332
rect 8018 19292 8024 19304
rect 7979 19264 8024 19292
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19292 9091 19295
rect 11146 19292 11152 19304
rect 9079 19264 10180 19292
rect 11107 19264 11152 19292
rect 9079 19261 9091 19264
rect 9033 19255 9091 19261
rect 9769 19227 9827 19233
rect 9769 19193 9781 19227
rect 9815 19224 9827 19227
rect 9858 19224 9864 19236
rect 9815 19196 9864 19224
rect 9815 19193 9827 19196
rect 9769 19187 9827 19193
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 8386 19156 8392 19168
rect 8347 19128 8392 19156
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 10152 19156 10180 19264
rect 11146 19252 11152 19264
rect 11204 19292 11210 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11204 19264 11529 19292
rect 11204 19252 11210 19264
rect 11517 19261 11529 19264
rect 11563 19292 11575 19295
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11563 19264 12265 19292
rect 11563 19261 11575 19264
rect 11517 19255 11575 19261
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 12253 19255 12311 19261
rect 14568 19264 14933 19292
rect 10502 19156 10508 19168
rect 10152 19128 10508 19156
rect 10502 19116 10508 19128
rect 10560 19156 10566 19168
rect 11238 19156 11244 19168
rect 10560 19128 11244 19156
rect 10560 19116 10566 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14568 19165 14596 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15930 19252 15936 19304
rect 15988 19292 15994 19304
rect 16592 19292 16620 19332
rect 17477 19329 17489 19332
rect 17523 19329 17535 19363
rect 17477 19323 17535 19329
rect 18046 19320 18052 19372
rect 18104 19360 18110 19372
rect 20548 19369 20576 19400
rect 21100 19369 21128 19468
rect 19133 19363 19191 19369
rect 19133 19360 19145 19363
rect 18104 19332 19145 19360
rect 18104 19320 18110 19332
rect 19133 19329 19145 19332
rect 19179 19329 19191 19363
rect 19133 19323 19191 19329
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 15988 19264 16620 19292
rect 17221 19295 17279 19301
rect 15988 19252 15994 19264
rect 17221 19261 17233 19295
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 13872 19128 13921 19156
rect 13872 19116 13878 19128
rect 13909 19125 13921 19128
rect 13955 19156 13967 19159
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 13955 19128 14565 19156
rect 13955 19125 13967 19128
rect 13909 19119 13967 19125
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 16298 19156 16304 19168
rect 16259 19128 16304 19156
rect 14553 19119 14611 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 17236 19156 17264 19255
rect 17954 19156 17960 19168
rect 16807 19128 17960 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17954 19116 17960 19128
rect 18012 19156 18018 19168
rect 18892 19156 18920 19255
rect 20254 19156 20260 19168
rect 18012 19128 18920 19156
rect 20215 19128 20260 19156
rect 18012 19116 18018 19128
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 20622 19116 20628 19168
rect 20680 19156 20686 19168
rect 20717 19159 20775 19165
rect 20717 19156 20729 19159
rect 20680 19128 20729 19156
rect 20680 19116 20686 19128
rect 20717 19125 20729 19128
rect 20763 19125 20775 19159
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 20717 19119 20775 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 11238 18952 11244 18964
rect 8076 18924 11100 18952
rect 11151 18924 11244 18952
rect 8076 18912 8082 18924
rect 11072 18884 11100 18924
rect 11238 18912 11244 18924
rect 11296 18952 11302 18964
rect 11698 18952 11704 18964
rect 11296 18924 11704 18952
rect 11296 18912 11302 18924
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 16298 18912 16304 18964
rect 16356 18952 16362 18964
rect 16356 18924 17724 18952
rect 16356 18912 16362 18924
rect 11882 18884 11888 18896
rect 11072 18856 11888 18884
rect 11882 18844 11888 18856
rect 11940 18844 11946 18896
rect 17586 18816 17592 18828
rect 17236 18788 17592 18816
rect 8205 18751 8263 18757
rect 8205 18717 8217 18751
rect 8251 18748 8263 18751
rect 8386 18748 8392 18760
rect 8251 18720 8392 18748
rect 8251 18717 8263 18720
rect 8205 18711 8263 18717
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 11146 18748 11152 18760
rect 9907 18720 11152 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 11146 18708 11152 18720
rect 11204 18748 11210 18760
rect 12897 18751 12955 18757
rect 11204 18720 12434 18748
rect 11204 18708 11210 18720
rect 9490 18640 9496 18692
rect 9548 18680 9554 18692
rect 10128 18683 10186 18689
rect 10128 18680 10140 18683
rect 9548 18652 10140 18680
rect 9548 18640 9554 18652
rect 10128 18649 10140 18652
rect 10174 18680 10186 18683
rect 10174 18652 11560 18680
rect 10174 18649 10186 18652
rect 10128 18643 10186 18649
rect 8386 18612 8392 18624
rect 8347 18584 8392 18612
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 11532 18621 11560 18652
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 9272 18584 9321 18612
rect 9272 18572 9278 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9309 18575 9367 18581
rect 11517 18615 11575 18621
rect 11517 18581 11529 18615
rect 11563 18581 11575 18615
rect 12406 18612 12434 18720
rect 12897 18717 12909 18751
rect 12943 18748 12955 18751
rect 13814 18748 13820 18760
rect 12943 18720 13820 18748
rect 12943 18717 12955 18720
rect 12897 18711 12955 18717
rect 12618 18640 12624 18692
rect 12676 18689 12682 18692
rect 12676 18680 12688 18689
rect 12676 18652 12721 18680
rect 12676 18643 12688 18652
rect 12676 18640 12682 18643
rect 12912 18612 12940 18711
rect 13814 18708 13820 18720
rect 13872 18748 13878 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13872 18720 14289 18748
rect 13872 18708 13878 18720
rect 14277 18717 14289 18720
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 14544 18751 14602 18757
rect 14544 18717 14556 18751
rect 14590 18748 14602 18751
rect 17236 18748 17264 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 17696 18816 17724 18924
rect 17696 18788 19380 18816
rect 14590 18720 17264 18748
rect 17313 18751 17371 18757
rect 14590 18717 14602 18720
rect 14544 18711 14602 18717
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 18690 18748 18696 18760
rect 17359 18720 17724 18748
rect 18651 18720 18696 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 17126 18689 17132 18692
rect 17068 18683 17132 18689
rect 17068 18680 17080 18683
rect 15672 18652 17080 18680
rect 13262 18612 13268 18624
rect 12406 18584 13268 18612
rect 11517 18575 11575 18581
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 15672 18621 15700 18652
rect 17068 18649 17080 18652
rect 17114 18649 17132 18683
rect 17068 18643 17132 18649
rect 17126 18640 17132 18643
rect 17184 18640 17190 18692
rect 15657 18615 15715 18621
rect 15657 18581 15669 18615
rect 15703 18581 15715 18615
rect 15930 18612 15936 18624
rect 15891 18584 15936 18612
rect 15657 18575 15715 18581
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 17696 18621 17724 18720
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19260 18680 19288 18711
rect 18340 18652 19288 18680
rect 19352 18680 19380 18788
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 22370 18748 22376 18760
rect 21131 18720 22376 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 22370 18708 22376 18720
rect 22428 18708 22434 18760
rect 19512 18683 19570 18689
rect 19512 18680 19524 18683
rect 19352 18652 19524 18680
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 17954 18612 17960 18624
rect 17727 18584 17960 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 17954 18572 17960 18584
rect 18012 18612 18018 18624
rect 18340 18621 18368 18652
rect 19512 18649 19524 18652
rect 19558 18680 19570 18683
rect 20346 18680 20352 18692
rect 19558 18652 20352 18680
rect 19558 18649 19570 18652
rect 19512 18643 19570 18649
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 18012 18584 18337 18612
rect 18012 18572 18018 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 18325 18575 18383 18581
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19150 18612 19156 18624
rect 18923 18584 19156 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 19944 18584 20637 18612
rect 19944 18572 19950 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 20772 18584 21281 18612
rect 20772 18572 20778 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 8849 18411 8907 18417
rect 8849 18408 8861 18411
rect 8628 18380 8861 18408
rect 8628 18368 8634 18380
rect 8849 18377 8861 18380
rect 8895 18377 8907 18411
rect 9214 18408 9220 18420
rect 9175 18380 9220 18408
rect 8849 18371 8907 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 11204 18380 11529 18408
rect 11204 18368 11210 18380
rect 11517 18377 11529 18380
rect 11563 18408 11575 18411
rect 11698 18408 11704 18420
rect 11563 18380 11704 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 11882 18368 11888 18420
rect 11940 18408 11946 18420
rect 12069 18411 12127 18417
rect 12069 18408 12081 18411
rect 11940 18380 12081 18408
rect 11940 18368 11946 18380
rect 12069 18377 12081 18380
rect 12115 18377 12127 18411
rect 12069 18371 12127 18377
rect 17310 18368 17316 18420
rect 17368 18408 17374 18420
rect 18969 18411 19027 18417
rect 18969 18408 18981 18411
rect 17368 18380 18981 18408
rect 17368 18368 17374 18380
rect 18969 18377 18981 18380
rect 19015 18377 19027 18411
rect 18969 18371 19027 18377
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 16942 18340 16948 18352
rect 8444 18312 16948 18340
rect 8444 18300 8450 18312
rect 16942 18300 16948 18312
rect 17000 18300 17006 18352
rect 13170 18232 13176 18284
rect 13228 18281 13234 18284
rect 13228 18272 13240 18281
rect 16045 18275 16103 18281
rect 13228 18244 13860 18272
rect 13228 18235 13240 18244
rect 13228 18232 13234 18235
rect 9306 18204 9312 18216
rect 9267 18176 9312 18204
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 9490 18204 9496 18216
rect 9451 18176 9496 18204
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 13449 18207 13507 18213
rect 13449 18173 13461 18207
rect 13495 18173 13507 18207
rect 13449 18167 13507 18173
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13464 18068 13492 18167
rect 13832 18136 13860 18244
rect 16045 18241 16057 18275
rect 16091 18272 16103 18275
rect 16758 18272 16764 18284
rect 16091 18244 16764 18272
rect 16091 18241 16103 18244
rect 16045 18235 16103 18241
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 17120 18275 17178 18281
rect 17120 18241 17132 18275
rect 17166 18272 17178 18275
rect 17494 18272 17500 18284
rect 17166 18244 17500 18272
rect 17166 18241 17178 18244
rect 17120 18235 17178 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 19150 18272 19156 18284
rect 19111 18244 19156 18272
rect 19150 18232 19156 18244
rect 19208 18232 19214 18284
rect 19429 18275 19487 18281
rect 19429 18241 19441 18275
rect 19475 18272 19487 18275
rect 19518 18272 19524 18284
rect 19475 18244 19524 18272
rect 19475 18241 19487 18244
rect 19429 18235 19487 18241
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 20254 18281 20260 18284
rect 20248 18272 20260 18281
rect 20215 18244 20260 18272
rect 20248 18235 20260 18244
rect 20254 18232 20260 18235
rect 20312 18232 20318 18284
rect 16298 18204 16304 18216
rect 16259 18176 16304 18204
rect 16298 18164 16304 18176
rect 16356 18204 16362 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 16356 18176 16865 18204
rect 16356 18164 16362 18176
rect 16853 18173 16865 18176
rect 16899 18173 16911 18207
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 16853 18167 16911 18173
rect 18524 18176 19993 18204
rect 14921 18139 14979 18145
rect 14921 18136 14933 18139
rect 13832 18108 14933 18136
rect 14921 18105 14933 18108
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 18524 18145 18552 18176
rect 19981 18173 19993 18176
rect 20027 18173 20039 18207
rect 19981 18167 20039 18173
rect 18509 18139 18567 18145
rect 18509 18136 18521 18139
rect 18012 18108 18521 18136
rect 18012 18096 18018 18108
rect 18509 18105 18521 18108
rect 18555 18105 18567 18139
rect 19610 18136 19616 18148
rect 19571 18108 19616 18136
rect 18509 18099 18567 18105
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 13725 18071 13783 18077
rect 13725 18068 13737 18071
rect 13320 18040 13737 18068
rect 13320 18028 13326 18040
rect 13725 18037 13737 18040
rect 13771 18068 13783 18071
rect 14553 18071 14611 18077
rect 14553 18068 14565 18071
rect 13771 18040 14565 18068
rect 13771 18037 13783 18040
rect 13725 18031 13783 18037
rect 14553 18037 14565 18040
rect 14599 18037 14611 18071
rect 14553 18031 14611 18037
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 18233 18071 18291 18077
rect 18233 18068 18245 18071
rect 18104 18040 18245 18068
rect 18104 18028 18110 18040
rect 18233 18037 18245 18040
rect 18279 18037 18291 18071
rect 18233 18031 18291 18037
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21542 18068 21548 18080
rect 21407 18040 21548 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 18874 17864 18880 17876
rect 18835 17836 18880 17864
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 20714 17864 20720 17876
rect 18984 17836 20720 17864
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 16485 17799 16543 17805
rect 16485 17796 16497 17799
rect 15620 17768 16497 17796
rect 15620 17756 15626 17768
rect 16485 17765 16497 17768
rect 16531 17765 16543 17799
rect 16485 17759 16543 17765
rect 18984 17728 19012 17836
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 17788 17700 19012 17728
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12906 17663 12964 17669
rect 12906 17660 12918 17663
rect 11940 17632 12918 17660
rect 11940 17620 11946 17632
rect 12906 17629 12918 17632
rect 12952 17629 12964 17663
rect 12906 17623 12964 17629
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17660 13231 17663
rect 17609 17663 17667 17669
rect 13219 17632 13308 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 13280 17536 13308 17632
rect 17609 17629 17621 17663
rect 17655 17660 17667 17663
rect 17788 17660 17816 17700
rect 17655 17632 17816 17660
rect 17865 17663 17923 17669
rect 17655 17629 17667 17632
rect 17609 17623 17667 17629
rect 17865 17629 17877 17663
rect 17911 17660 17923 17663
rect 17954 17660 17960 17672
rect 17911 17632 17960 17660
rect 17911 17629 17923 17632
rect 17865 17623 17923 17629
rect 17954 17620 17960 17632
rect 18012 17660 18018 17672
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 18012 17632 18153 17660
rect 18012 17620 18018 17632
rect 18141 17629 18153 17632
rect 18187 17629 18199 17663
rect 18141 17623 18199 17629
rect 18598 17620 18604 17672
rect 18656 17660 18662 17672
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 18656 17632 18705 17660
rect 18656 17620 18662 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 20625 17663 20683 17669
rect 20625 17660 20637 17663
rect 19300 17632 20637 17660
rect 19300 17620 19306 17632
rect 20625 17629 20637 17632
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17660 21143 17663
rect 21174 17660 21180 17672
rect 21131 17632 21180 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 19886 17552 19892 17604
rect 19944 17592 19950 17604
rect 20358 17595 20416 17601
rect 20358 17592 20370 17595
rect 19944 17564 20370 17592
rect 19944 17552 19950 17564
rect 20358 17561 20370 17564
rect 20404 17561 20416 17595
rect 20358 17555 20416 17561
rect 11790 17524 11796 17536
rect 11751 17496 11796 17524
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13320 17496 13461 17524
rect 13320 17484 13326 17496
rect 13449 17493 13461 17496
rect 13495 17524 13507 17527
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 13495 17496 15025 17524
rect 13495 17493 13507 17496
rect 13449 17487 13507 17493
rect 15013 17493 15025 17496
rect 15059 17524 15071 17527
rect 15381 17527 15439 17533
rect 15381 17524 15393 17527
rect 15059 17496 15393 17524
rect 15059 17493 15071 17496
rect 15013 17487 15071 17493
rect 15381 17493 15393 17496
rect 15427 17524 15439 17527
rect 15749 17527 15807 17533
rect 15749 17524 15761 17527
rect 15427 17496 15761 17524
rect 15427 17493 15439 17496
rect 15381 17487 15439 17493
rect 15749 17493 15761 17496
rect 15795 17524 15807 17527
rect 15838 17524 15844 17536
rect 15795 17496 15844 17524
rect 15795 17493 15807 17496
rect 15749 17487 15807 17493
rect 15838 17484 15844 17496
rect 15896 17524 15902 17536
rect 16117 17527 16175 17533
rect 16117 17524 16129 17527
rect 15896 17496 16129 17524
rect 15896 17484 15902 17496
rect 16117 17493 16129 17496
rect 16163 17524 16175 17527
rect 16298 17524 16304 17536
rect 16163 17496 16304 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 19245 17527 19303 17533
rect 19245 17493 19257 17527
rect 19291 17524 19303 17527
rect 19702 17524 19708 17536
rect 19291 17496 19708 17524
rect 19291 17493 19303 17496
rect 19245 17487 19303 17493
rect 19702 17484 19708 17496
rect 19760 17524 19766 17536
rect 20254 17524 20260 17536
rect 19760 17496 20260 17524
rect 19760 17484 19766 17496
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 20530 17484 20536 17536
rect 20588 17524 20594 17536
rect 21269 17527 21327 17533
rect 21269 17524 21281 17527
rect 20588 17496 21281 17524
rect 20588 17484 20594 17496
rect 21269 17493 21281 17496
rect 21315 17493 21327 17527
rect 21269 17487 21327 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 11698 17320 11704 17332
rect 11659 17292 11704 17320
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 11716 17184 11744 17280
rect 15838 17212 15844 17264
rect 15896 17252 15902 17264
rect 16669 17255 16727 17261
rect 16669 17252 16681 17255
rect 15896 17224 16681 17252
rect 15896 17212 15902 17224
rect 16669 17221 16681 17224
rect 16715 17221 16727 17255
rect 16669 17215 16727 17221
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 20438 17252 20444 17264
rect 18012 17224 18644 17252
rect 18012 17212 18018 17224
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11716 17156 12081 17184
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12336 17187 12394 17193
rect 12336 17153 12348 17187
rect 12382 17184 12394 17187
rect 13722 17184 13728 17196
rect 12382 17156 13728 17184
rect 12382 17153 12394 17156
rect 12336 17147 12394 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 15188 17187 15246 17193
rect 15188 17153 15200 17187
rect 15234 17184 15246 17187
rect 15562 17184 15568 17196
rect 15234 17156 15568 17184
rect 15234 17153 15246 17156
rect 15188 17147 15246 17153
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 18345 17187 18403 17193
rect 18345 17153 18357 17187
rect 18391 17184 18403 17187
rect 18506 17184 18512 17196
rect 18391 17156 18512 17184
rect 18391 17153 18403 17156
rect 18345 17147 18403 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18616 17193 18644 17224
rect 19168 17224 20444 17252
rect 19168 17193 19196 17224
rect 20438 17212 20444 17224
rect 20496 17212 20502 17264
rect 19702 17193 19708 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 19696 17147 19708 17193
rect 19760 17184 19766 17196
rect 21082 17184 21088 17196
rect 19760 17156 19796 17184
rect 21043 17156 21088 17184
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 13740 17088 14933 17116
rect 13262 17008 13268 17060
rect 13320 17048 13326 17060
rect 13740 17057 13768 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 18616 17116 18644 17147
rect 19702 17144 19708 17147
rect 19760 17144 19766 17156
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 19242 17116 19248 17128
rect 18616 17088 19248 17116
rect 14921 17079 14979 17085
rect 19242 17076 19248 17088
rect 19300 17116 19306 17128
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 19300 17088 19441 17116
rect 19300 17076 19306 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 13320 17020 13737 17048
rect 13320 17008 13326 17020
rect 13725 17017 13737 17020
rect 13771 17017 13783 17051
rect 13725 17011 13783 17017
rect 16301 17051 16359 17057
rect 16301 17017 16313 17051
rect 16347 17048 16359 17051
rect 17310 17048 17316 17060
rect 16347 17020 17316 17048
rect 16347 17017 16359 17020
rect 16301 17011 16359 17017
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 18966 17048 18972 17060
rect 18927 17020 18972 17048
rect 18966 17008 18972 17020
rect 19024 17008 19030 17060
rect 20622 17008 20628 17060
rect 20680 17048 20686 17060
rect 21269 17051 21327 17057
rect 21269 17048 21281 17051
rect 20680 17020 21281 17048
rect 20680 17008 20686 17020
rect 21269 17017 21281 17020
rect 21315 17017 21327 17051
rect 21269 17011 21327 17017
rect 13449 16983 13507 16989
rect 13449 16949 13461 16983
rect 13495 16980 13507 16983
rect 14550 16980 14556 16992
rect 13495 16952 14556 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 17221 16983 17279 16989
rect 17221 16949 17233 16983
rect 17267 16980 17279 16983
rect 17678 16980 17684 16992
rect 17267 16952 17684 16980
rect 17267 16949 17279 16952
rect 17221 16943 17279 16949
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 20809 16983 20867 16989
rect 20809 16980 20821 16983
rect 20772 16952 20821 16980
rect 20772 16940 20778 16952
rect 20809 16949 20821 16952
rect 20855 16980 20867 16983
rect 22738 16980 22744 16992
rect 20855 16952 22744 16980
rect 20855 16949 20867 16952
rect 20809 16943 20867 16949
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 10502 16776 10508 16788
rect 10463 16748 10508 16776
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 11756 16748 11928 16776
rect 11756 16736 11762 16748
rect 9953 16711 10011 16717
rect 9953 16708 9965 16711
rect 9416 16680 9965 16708
rect 9416 16652 9444 16680
rect 9953 16677 9965 16680
rect 9999 16677 10011 16711
rect 9953 16671 10011 16677
rect 9398 16640 9404 16652
rect 9311 16612 9404 16640
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16640 9643 16643
rect 9858 16640 9864 16652
rect 9631 16612 9864 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 11900 16649 11928 16748
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 18782 16776 18788 16788
rect 18564 16748 18788 16776
rect 18564 16736 18570 16748
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 11931 16612 12173 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12161 16609 12173 16612
rect 12207 16609 12219 16643
rect 12161 16603 12219 16609
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 14277 16643 14335 16649
rect 14277 16640 14289 16643
rect 13320 16612 14289 16640
rect 13320 16600 13326 16612
rect 14277 16609 14289 16612
rect 14323 16609 14335 16643
rect 14277 16603 14335 16609
rect 11629 16575 11687 16581
rect 11629 16541 11641 16575
rect 11675 16572 11687 16575
rect 11790 16572 11796 16584
rect 11675 16544 11796 16572
rect 11675 16541 11687 16544
rect 11629 16535 11687 16541
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 15933 16575 15991 16581
rect 15933 16572 15945 16575
rect 15896 16544 15945 16572
rect 15896 16532 15902 16544
rect 15933 16541 15945 16544
rect 15979 16572 15991 16575
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 15979 16544 17601 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 17589 16541 17601 16544
rect 17635 16572 17647 16575
rect 17954 16572 17960 16584
rect 17635 16544 17960 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17954 16532 17960 16544
rect 18012 16572 18018 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18012 16544 18337 16572
rect 18012 16532 18018 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 14550 16513 14556 16516
rect 9309 16507 9367 16513
rect 9309 16504 9321 16507
rect 8496 16476 9321 16504
rect 8496 16448 8524 16476
rect 9309 16473 9321 16476
rect 9355 16473 9367 16507
rect 12406 16507 12464 16513
rect 12406 16504 12418 16507
rect 9309 16467 9367 16473
rect 11716 16476 12418 16504
rect 8478 16436 8484 16448
rect 8439 16408 8484 16436
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8720 16408 8953 16436
rect 8720 16396 8726 16408
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11716 16436 11744 16476
rect 12406 16473 12418 16476
rect 12452 16473 12464 16507
rect 14544 16504 14556 16513
rect 14511 16476 14556 16504
rect 12406 16467 12464 16473
rect 14544 16467 14556 16476
rect 14550 16464 14556 16467
rect 14608 16464 14614 16516
rect 16206 16513 16212 16516
rect 16200 16504 16212 16513
rect 15672 16476 16212 16504
rect 11020 16408 11744 16436
rect 13541 16439 13599 16445
rect 11020 16396 11026 16408
rect 13541 16405 13553 16439
rect 13587 16436 13599 16439
rect 13722 16436 13728 16448
rect 13587 16408 13728 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 15672 16445 15700 16476
rect 16200 16467 16212 16476
rect 16206 16464 16212 16467
rect 16264 16464 16270 16516
rect 17862 16464 17868 16516
rect 17920 16504 17926 16516
rect 18708 16504 18736 16535
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 19300 16544 20637 16572
rect 19300 16532 19306 16544
rect 20625 16541 20637 16544
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16572 21143 16575
rect 22186 16572 22192 16584
rect 21131 16544 22192 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 19518 16504 19524 16516
rect 17920 16476 18736 16504
rect 18892 16476 19524 16504
rect 17920 16464 17926 16476
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16405 15715 16439
rect 15657 16399 15715 16405
rect 17313 16439 17371 16445
rect 17313 16405 17325 16439
rect 17359 16436 17371 16439
rect 17494 16436 17500 16448
rect 17359 16408 17500 16436
rect 17359 16405 17371 16408
rect 17313 16399 17371 16405
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 18892 16445 18920 16476
rect 19518 16464 19524 16476
rect 19576 16464 19582 16516
rect 20380 16507 20438 16513
rect 20380 16473 20392 16507
rect 20426 16504 20438 16507
rect 20806 16504 20812 16516
rect 20426 16476 20812 16504
rect 20426 16473 20438 16476
rect 20380 16467 20438 16473
rect 20806 16464 20812 16476
rect 20864 16504 20870 16516
rect 22094 16504 22100 16516
rect 20864 16476 22100 16504
rect 20864 16464 20870 16476
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 18877 16439 18935 16445
rect 18877 16405 18889 16439
rect 18923 16405 18935 16439
rect 18877 16399 18935 16405
rect 19245 16439 19303 16445
rect 19245 16405 19257 16439
rect 19291 16436 19303 16439
rect 20070 16436 20076 16448
rect 19291 16408 20076 16436
rect 19291 16405 19303 16408
rect 19245 16399 19303 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 21266 16436 21272 16448
rect 21227 16408 21272 16436
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 15838 16232 15844 16244
rect 15799 16204 15844 16232
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 19150 16192 19156 16244
rect 19208 16232 19214 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 19208 16204 19441 16232
rect 19208 16192 19214 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 20714 16164 20720 16176
rect 19628 16136 20720 16164
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 12630 16099 12688 16105
rect 12630 16096 12642 16099
rect 9640 16068 12642 16096
rect 9640 16056 9646 16068
rect 12630 16065 12642 16068
rect 12676 16065 12688 16099
rect 12630 16059 12688 16065
rect 17793 16099 17851 16105
rect 17793 16065 17805 16099
rect 17839 16096 17851 16099
rect 17954 16096 17960 16108
rect 17839 16068 17960 16096
rect 17839 16065 17851 16068
rect 17793 16059 17851 16065
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 19628 16105 19656 16136
rect 20714 16124 20720 16136
rect 20772 16124 20778 16176
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 20145 16099 20203 16105
rect 20145 16096 20157 16099
rect 19852 16068 20157 16096
rect 19852 16056 19858 16068
rect 20145 16065 20157 16068
rect 20191 16065 20203 16099
rect 20145 16059 20203 16065
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 16028 12955 16031
rect 18046 16028 18052 16040
rect 12943 16000 13308 16028
rect 18007 16000 18052 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 13280 15904 13308 16000
rect 18046 15988 18052 16000
rect 18104 16028 18110 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18104 16000 18337 16028
rect 18104 15988 18110 16000
rect 18325 15997 18337 16000
rect 18371 16028 18383 16031
rect 18969 16031 19027 16037
rect 18969 16028 18981 16031
rect 18371 16000 18981 16028
rect 18371 15997 18383 16000
rect 18325 15991 18383 15997
rect 18969 15997 18981 16000
rect 19015 16028 19027 16031
rect 19242 16028 19248 16040
rect 19015 16000 19248 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 19242 15988 19248 16000
rect 19300 16028 19306 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19300 16000 19901 16028
rect 19300 15988 19306 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10962 15892 10968 15904
rect 9916 15864 10968 15892
rect 9916 15852 9922 15864
rect 10962 15852 10968 15864
rect 11020 15892 11026 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11020 15864 11529 15892
rect 11020 15852 11026 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 13262 15892 13268 15904
rect 13223 15864 13268 15892
rect 11517 15855 11575 15861
rect 13262 15852 13268 15864
rect 13320 15892 13326 15904
rect 13633 15895 13691 15901
rect 13633 15892 13645 15895
rect 13320 15864 13645 15892
rect 13320 15852 13326 15864
rect 13633 15861 13645 15864
rect 13679 15861 13691 15895
rect 13633 15855 13691 15861
rect 16669 15895 16727 15901
rect 16669 15861 16681 15895
rect 16715 15892 16727 15895
rect 16942 15892 16948 15904
rect 16715 15864 16948 15892
rect 16715 15861 16727 15864
rect 16669 15855 16727 15861
rect 16942 15852 16948 15864
rect 17000 15892 17006 15904
rect 17402 15892 17408 15904
rect 17000 15864 17408 15892
rect 17000 15852 17006 15864
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 20990 15852 20996 15904
rect 21048 15892 21054 15904
rect 21269 15895 21327 15901
rect 21269 15892 21281 15895
rect 21048 15864 21281 15892
rect 21048 15852 21054 15864
rect 21269 15861 21281 15864
rect 21315 15861 21327 15895
rect 21269 15855 21327 15861
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 21634 15688 21640 15700
rect 19720 15660 21640 15688
rect 15838 15552 15844 15564
rect 15799 15524 15844 15552
rect 15838 15512 15844 15524
rect 15896 15552 15902 15564
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15896 15524 16129 15552
rect 15896 15512 15902 15524
rect 16117 15521 16129 15524
rect 16163 15552 16175 15555
rect 16298 15552 16304 15564
rect 16163 15524 16304 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16298 15512 16304 15524
rect 16356 15552 16362 15564
rect 16485 15555 16543 15561
rect 16485 15552 16497 15555
rect 16356 15524 16497 15552
rect 16356 15512 16362 15524
rect 16485 15521 16497 15524
rect 16531 15552 16543 15555
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 16531 15524 17049 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 17037 15521 17049 15524
rect 17083 15552 17095 15555
rect 17405 15555 17463 15561
rect 17405 15552 17417 15555
rect 17083 15524 17417 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 17405 15521 17417 15524
rect 17451 15552 17463 15555
rect 17773 15555 17831 15561
rect 17773 15552 17785 15555
rect 17451 15524 17785 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 17773 15521 17785 15524
rect 17819 15552 17831 15555
rect 18046 15552 18052 15564
rect 17819 15524 18052 15552
rect 17819 15521 17831 15524
rect 17773 15515 17831 15521
rect 18046 15512 18052 15524
rect 18104 15552 18110 15564
rect 18141 15555 18199 15561
rect 18141 15552 18153 15555
rect 18104 15524 18153 15552
rect 18104 15512 18110 15524
rect 18141 15521 18153 15524
rect 18187 15552 18199 15555
rect 18785 15555 18843 15561
rect 18785 15552 18797 15555
rect 18187 15524 18797 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18785 15521 18797 15524
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 19720 15493 19748 15660
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15484 12495 15487
rect 19705 15487 19763 15493
rect 12483 15456 12848 15484
rect 12483 15453 12495 15456
rect 12437 15447 12495 15453
rect 12066 15376 12072 15428
rect 12124 15416 12130 15428
rect 12170 15419 12228 15425
rect 12170 15416 12182 15419
rect 12124 15388 12182 15416
rect 12124 15376 12130 15388
rect 12170 15385 12182 15388
rect 12216 15385 12228 15419
rect 12170 15379 12228 15385
rect 9582 15308 9588 15360
rect 9640 15348 9646 15360
rect 12820 15357 12848 15456
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 20680 15456 21373 15484
rect 20680 15444 20686 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 15596 15419 15654 15425
rect 15596 15385 15608 15419
rect 15642 15416 15654 15419
rect 18230 15416 18236 15428
rect 15642 15388 18236 15416
rect 15642 15385 15654 15388
rect 15596 15379 15654 15385
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 21116 15419 21174 15425
rect 21116 15385 21128 15419
rect 21162 15416 21174 15419
rect 21162 15388 21404 15416
rect 21162 15385 21174 15388
rect 21116 15379 21174 15385
rect 21376 15360 21404 15388
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 9640 15320 11069 15348
rect 9640 15308 9646 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 12805 15351 12863 15357
rect 12805 15317 12817 15351
rect 12851 15348 12863 15351
rect 13262 15348 13268 15360
rect 12851 15320 13268 15348
rect 12851 15317 12863 15320
rect 12805 15311 12863 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 14461 15351 14519 15357
rect 14461 15317 14473 15351
rect 14507 15348 14519 15351
rect 14826 15348 14832 15360
rect 14507 15320 14832 15348
rect 14507 15317 14519 15320
rect 14461 15311 14519 15317
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 19242 15308 19248 15360
rect 19300 15348 19306 15360
rect 19521 15351 19579 15357
rect 19521 15348 19533 15351
rect 19300 15320 19533 15348
rect 19300 15308 19306 15320
rect 19521 15317 19533 15320
rect 19567 15317 19579 15351
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19521 15311 19579 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 21358 15308 21364 15360
rect 21416 15308 21422 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 16298 15144 16304 15156
rect 16259 15116 16304 15144
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 18322 15144 18328 15156
rect 17880 15116 18328 15144
rect 17793 15079 17851 15085
rect 17793 15045 17805 15079
rect 17839 15076 17851 15079
rect 17880 15076 17908 15116
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 20622 15076 20628 15088
rect 17839 15048 17908 15076
rect 18064 15048 20628 15076
rect 17839 15045 17851 15048
rect 17793 15039 17851 15045
rect 18064 15020 18092 15048
rect 13009 15011 13067 15017
rect 13009 14977 13021 15011
rect 13055 15008 13067 15011
rect 13814 15008 13820 15020
rect 13055 14980 13820 15008
rect 13055 14977 13067 14980
rect 13009 14971 13067 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14826 15017 14832 15020
rect 14820 15008 14832 15017
rect 14787 14980 14832 15008
rect 14820 14971 14832 14980
rect 14826 14968 14832 14971
rect 14884 14968 14890 15020
rect 18046 15008 18052 15020
rect 18007 14980 18052 15008
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 19720 15017 19748 15048
rect 20622 15036 20628 15048
rect 20680 15076 20686 15088
rect 20680 15048 21404 15076
rect 20680 15036 20686 15048
rect 19449 15011 19507 15017
rect 19449 14977 19461 15011
rect 19495 15008 19507 15011
rect 19705 15011 19763 15017
rect 19495 14980 19656 15008
rect 19495 14977 19507 14980
rect 19449 14971 19507 14977
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 13320 14912 14565 14940
rect 13320 14900 13326 14912
rect 13648 14816 13676 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 19628 14940 19656 14980
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 20806 15008 20812 15020
rect 19705 14971 19763 14977
rect 19812 14980 20812 15008
rect 19812 14940 19840 14980
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 21376 15017 21404 15048
rect 21105 15011 21163 15017
rect 21105 14977 21117 15011
rect 21151 15008 21163 15011
rect 21361 15011 21419 15017
rect 21151 14980 21312 15008
rect 21151 14977 21163 14980
rect 21105 14971 21163 14977
rect 19628 14912 19840 14940
rect 21284 14940 21312 14980
rect 21361 14977 21373 15011
rect 21407 14977 21419 15011
rect 21361 14971 21419 14977
rect 21450 14940 21456 14952
rect 21284 14912 21456 14940
rect 14553 14903 14611 14909
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 15933 14875 15991 14881
rect 15933 14841 15945 14875
rect 15979 14872 15991 14875
rect 15979 14844 17172 14872
rect 15979 14841 15991 14844
rect 15933 14835 15991 14841
rect 11885 14807 11943 14813
rect 11885 14773 11897 14807
rect 11931 14804 11943 14807
rect 12066 14804 12072 14816
rect 11931 14776 12072 14804
rect 11931 14773 11943 14776
rect 11885 14767 11943 14773
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 13630 14804 13636 14816
rect 13591 14776 13636 14804
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 16666 14804 16672 14816
rect 16627 14776 16672 14804
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17144 14804 17172 14844
rect 18138 14804 18144 14816
rect 17144 14776 18144 14804
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 18288 14776 18337 14804
rect 18288 14764 18294 14776
rect 18325 14773 18337 14776
rect 18371 14804 18383 14807
rect 18966 14804 18972 14816
rect 18371 14776 18972 14804
rect 18371 14773 18383 14776
rect 18325 14767 18383 14773
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19794 14764 19800 14816
rect 19852 14804 19858 14816
rect 19981 14807 20039 14813
rect 19981 14804 19993 14807
rect 19852 14776 19993 14804
rect 19852 14764 19858 14776
rect 19981 14773 19993 14776
rect 20027 14773 20039 14807
rect 19981 14767 20039 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 18046 14600 18052 14612
rect 14884 14572 18052 14600
rect 14884 14560 14890 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19518 14600 19524 14612
rect 19479 14572 19524 14600
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 16117 14535 16175 14541
rect 16117 14501 16129 14535
rect 16163 14501 16175 14535
rect 16117 14495 16175 14501
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 12032 14368 12081 14396
rect 12032 14356 12038 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13688 14368 13737 14396
rect 13688 14356 13694 14368
rect 13725 14365 13737 14368
rect 13771 14396 13783 14399
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13771 14368 14105 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14139 14368 14473 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 15930 14396 15936 14408
rect 14461 14359 14519 14365
rect 14660 14368 15936 14396
rect 11824 14331 11882 14337
rect 11824 14297 11836 14331
rect 11870 14328 11882 14331
rect 13480 14331 13538 14337
rect 11870 14300 12388 14328
rect 11870 14297 11882 14300
rect 11824 14291 11882 14297
rect 10689 14263 10747 14269
rect 10689 14229 10701 14263
rect 10735 14260 10747 14263
rect 11698 14260 11704 14272
rect 10735 14232 11704 14260
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12360 14269 12388 14300
rect 13480 14297 13492 14331
rect 13526 14328 13538 14331
rect 14660 14328 14688 14368
rect 15930 14356 15936 14368
rect 15988 14396 15994 14408
rect 16132 14396 16160 14495
rect 15988 14368 16160 14396
rect 15988 14356 15994 14368
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 16356 14368 17509 14396
rect 16356 14356 16362 14368
rect 17497 14365 17509 14368
rect 17543 14396 17555 14399
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17543 14368 17785 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 17773 14365 17785 14368
rect 17819 14396 17831 14399
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 17819 14368 18337 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18325 14365 18337 14368
rect 18371 14396 18383 14399
rect 18506 14396 18512 14408
rect 18371 14368 18512 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18506 14356 18512 14368
rect 18564 14396 18570 14408
rect 18785 14399 18843 14405
rect 18785 14396 18797 14399
rect 18564 14368 18797 14396
rect 18564 14356 18570 14368
rect 18785 14365 18797 14368
rect 18831 14365 18843 14399
rect 19702 14396 19708 14408
rect 19663 14368 19708 14396
rect 18785 14359 18843 14365
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 20622 14356 20628 14408
rect 20680 14396 20686 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20680 14368 21373 14396
rect 20680 14356 20686 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 13526 14300 14688 14328
rect 14728 14331 14786 14337
rect 13526 14297 13538 14300
rect 13480 14291 13538 14297
rect 14728 14297 14740 14331
rect 14774 14328 14786 14331
rect 16942 14328 16948 14340
rect 14774 14300 16948 14328
rect 14774 14297 14786 14300
rect 14728 14291 14786 14297
rect 16942 14288 16948 14300
rect 17000 14288 17006 14340
rect 17218 14288 17224 14340
rect 17276 14337 17282 14340
rect 17276 14331 17299 14337
rect 17287 14297 17299 14331
rect 17276 14291 17299 14297
rect 17276 14288 17282 14291
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 21094 14331 21152 14337
rect 21094 14328 21106 14331
rect 21048 14300 21106 14328
rect 21048 14288 21054 14300
rect 21094 14297 21106 14300
rect 21140 14297 21152 14331
rect 21094 14291 21152 14297
rect 12345 14263 12403 14269
rect 12345 14229 12357 14263
rect 12391 14260 12403 14263
rect 12894 14260 12900 14272
rect 12391 14232 12900 14260
rect 12391 14229 12403 14232
rect 12345 14223 12403 14229
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 15841 14263 15899 14269
rect 15841 14229 15853 14263
rect 15887 14260 15899 14263
rect 18322 14260 18328 14272
rect 15887 14232 18328 14260
rect 15887 14229 15899 14232
rect 15841 14223 15899 14229
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 19981 14263 20039 14269
rect 19981 14229 19993 14263
rect 20027 14260 20039 14263
rect 20806 14260 20812 14272
rect 20027 14232 20812 14260
rect 20027 14229 20039 14232
rect 19981 14223 20039 14229
rect 20806 14220 20812 14232
rect 20864 14260 20870 14272
rect 22646 14260 22652 14272
rect 20864 14232 22652 14260
rect 20864 14220 20870 14232
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 8665 14059 8723 14065
rect 8665 14025 8677 14059
rect 8711 14056 8723 14059
rect 10042 14056 10048 14068
rect 8711 14028 10048 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 13357 14059 13415 14065
rect 13357 14025 13369 14059
rect 13403 14056 13415 14059
rect 13814 14056 13820 14068
rect 13403 14028 13820 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17678 14056 17684 14068
rect 17000 14028 17684 14056
rect 17000 14016 17006 14028
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 18233 14059 18291 14065
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 18414 14056 18420 14068
rect 18279 14028 18420 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 18414 14016 18420 14028
rect 18472 14056 18478 14068
rect 19610 14056 19616 14068
rect 18472 14028 19616 14056
rect 18472 14016 18478 14028
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 19889 14059 19947 14065
rect 19889 14025 19901 14059
rect 19935 14056 19947 14059
rect 20714 14056 20720 14068
rect 19935 14028 20576 14056
rect 20675 14028 20720 14056
rect 19935 14025 19947 14028
rect 19889 14019 19947 14025
rect 8205 13991 8263 13997
rect 8205 13957 8217 13991
rect 8251 13988 8263 13991
rect 9033 13991 9091 13997
rect 9033 13988 9045 13991
rect 8251 13960 9045 13988
rect 8251 13957 8263 13960
rect 8205 13951 8263 13957
rect 9033 13957 9045 13960
rect 9079 13988 9091 13991
rect 9398 13988 9404 14000
rect 9079 13960 9404 13988
rect 9079 13957 9091 13960
rect 9033 13951 9091 13957
rect 9398 13948 9404 13960
rect 9456 13988 9462 14000
rect 15746 13988 15752 14000
rect 9456 13960 15752 13988
rect 9456 13948 9462 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 17120 13991 17178 13997
rect 17120 13957 17132 13991
rect 17166 13988 17178 13991
rect 17218 13988 17224 14000
rect 17166 13960 17224 13988
rect 17166 13957 17178 13960
rect 17120 13951 17178 13957
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 18776 13991 18834 13997
rect 18776 13957 18788 13991
rect 18822 13988 18834 13991
rect 18874 13988 18880 14000
rect 18822 13960 18880 13988
rect 18822 13957 18834 13960
rect 18776 13951 18834 13957
rect 18874 13948 18880 13960
rect 18932 13988 18938 14000
rect 19978 13988 19984 14000
rect 18932 13960 19984 13988
rect 18932 13948 18938 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20548 13988 20576 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 21450 13988 21456 14000
rect 20548 13960 21456 13988
rect 21450 13948 21456 13960
rect 21508 13988 21514 14000
rect 22278 13988 22284 14000
rect 21508 13960 22284 13988
rect 21508 13948 21514 13960
rect 22278 13948 22284 13960
rect 22336 13948 22342 14000
rect 8294 13920 8300 13932
rect 8255 13892 8300 13920
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 12244 13923 12302 13929
rect 12244 13889 12256 13923
rect 12290 13920 12302 13923
rect 12802 13920 12808 13932
rect 12290 13892 12808 13920
rect 12290 13889 12302 13892
rect 12244 13883 12302 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16356 13892 16865 13920
rect 16356 13880 16362 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 18506 13920 18512 13932
rect 18467 13892 18512 13920
rect 16853 13883 16911 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 20530 13920 20536 13932
rect 20491 13892 20536 13920
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20990 13880 20996 13932
rect 21048 13920 21054 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 21048 13892 21097 13920
rect 21048 13880 21054 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 8113 13855 8171 13861
rect 8113 13821 8125 13855
rect 8159 13821 8171 13855
rect 11974 13852 11980 13864
rect 8113 13815 8171 13821
rect 11624 13824 11980 13852
rect 8128 13784 8156 13815
rect 9582 13784 9588 13796
rect 8128 13756 9588 13784
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11624 13725 11652 13824
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 16022 13852 16028 13864
rect 15983 13824 16028 13852
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 21450 13852 21456 13864
rect 20680 13824 21456 13852
rect 20680 13812 20686 13824
rect 21450 13812 21456 13824
rect 21508 13812 21514 13864
rect 11609 13719 11667 13725
rect 11609 13716 11621 13719
rect 11204 13688 11621 13716
rect 11204 13676 11210 13688
rect 11609 13685 11621 13688
rect 11655 13685 11667 13719
rect 13630 13716 13636 13728
rect 13591 13688 13636 13716
rect 11609 13679 11667 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 17494 13716 17500 13728
rect 17184 13688 17500 13716
rect 17184 13676 17190 13688
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20165 13719 20223 13725
rect 20165 13716 20177 13719
rect 20036 13688 20177 13716
rect 20036 13676 20042 13688
rect 20165 13685 20177 13688
rect 20211 13685 20223 13719
rect 21266 13716 21272 13728
rect 21227 13688 21272 13716
rect 20165 13679 20223 13685
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 21358 13512 21364 13524
rect 21319 13484 21364 13512
rect 21358 13472 21364 13484
rect 21416 13512 21422 13524
rect 22554 13512 22560 13524
rect 21416 13484 22560 13512
rect 21416 13472 21422 13484
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 11146 13376 11152 13388
rect 11107 13348 11152 13376
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14608 13348 15669 13376
rect 14608 13336 14614 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 18417 13379 18475 13385
rect 18417 13345 18429 13379
rect 18463 13376 18475 13379
rect 18506 13376 18512 13388
rect 18463 13348 18512 13376
rect 18463 13345 18475 13348
rect 18417 13339 18475 13345
rect 18506 13336 18512 13348
rect 18564 13376 18570 13388
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 18564 13348 18705 13376
rect 18564 13336 18570 13348
rect 18693 13345 18705 13348
rect 18739 13376 18751 13379
rect 19978 13376 19984 13388
rect 18739 13348 19984 13376
rect 18739 13345 18751 13348
rect 18693 13339 18751 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 11164 13308 11192 13336
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 11164 13280 12817 13308
rect 12805 13277 12817 13280
rect 12851 13308 12863 13311
rect 13630 13308 13636 13320
rect 12851 13280 13636 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16022 13308 16028 13320
rect 15979 13280 16028 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 16172 13280 19533 13308
rect 16172 13268 16178 13280
rect 19521 13277 19533 13280
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 20070 13268 20076 13320
rect 20128 13308 20134 13320
rect 20237 13311 20295 13317
rect 20237 13308 20249 13311
rect 20128 13280 20249 13308
rect 20128 13268 20134 13280
rect 20237 13277 20249 13280
rect 20283 13308 20295 13311
rect 20283 13280 20392 13308
rect 20283 13277 20295 13280
rect 20237 13271 20295 13277
rect 20364 13252 20392 13280
rect 11416 13243 11474 13249
rect 11416 13209 11428 13243
rect 11462 13240 11474 13243
rect 11698 13240 11704 13252
rect 11462 13212 11704 13240
rect 11462 13209 11474 13212
rect 11416 13203 11474 13209
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 17954 13240 17960 13252
rect 16316 13212 17960 13240
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12802 13172 12808 13184
rect 12575 13144 12808 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 15841 13175 15899 13181
rect 15841 13141 15853 13175
rect 15887 13172 15899 13175
rect 16206 13172 16212 13184
rect 15887 13144 16212 13172
rect 15887 13141 15899 13144
rect 15841 13135 15899 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 16316 13181 16344 13212
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 18138 13200 18144 13252
rect 18196 13249 18202 13252
rect 18196 13240 18208 13249
rect 18196 13212 18241 13240
rect 18196 13203 18208 13212
rect 18196 13200 18202 13203
rect 20346 13200 20352 13252
rect 20404 13200 20410 13252
rect 16301 13175 16359 13181
rect 16301 13141 16313 13175
rect 16347 13141 16359 13175
rect 16301 13135 16359 13141
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 16577 13175 16635 13181
rect 16577 13172 16589 13175
rect 16448 13144 16589 13172
rect 16448 13132 16454 13144
rect 16577 13141 16589 13144
rect 16623 13141 16635 13175
rect 16577 13135 16635 13141
rect 17037 13175 17095 13181
rect 17037 13141 17049 13175
rect 17083 13172 17095 13175
rect 17218 13172 17224 13184
rect 17083 13144 17224 13172
rect 17083 13141 17095 13144
rect 17037 13135 17095 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 19705 13175 19763 13181
rect 19705 13141 19717 13175
rect 19751 13172 19763 13175
rect 20714 13172 20720 13184
rect 19751 13144 20720 13172
rect 19751 13141 19763 13144
rect 19705 13135 19763 13141
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 15473 12971 15531 12977
rect 15473 12937 15485 12971
rect 15519 12968 15531 12971
rect 16114 12968 16120 12980
rect 15519 12940 16120 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 18690 12968 18696 12980
rect 18651 12940 18696 12968
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 20809 12971 20867 12977
rect 20809 12937 20821 12971
rect 20855 12968 20867 12971
rect 21082 12968 21088 12980
rect 20855 12940 21088 12968
rect 20855 12937 20867 12940
rect 20809 12931 20867 12937
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 18966 12900 18972 12912
rect 17543 12872 18972 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15151 12804 15761 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12832 17463 12835
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 17451 12804 18061 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 18049 12801 18061 12804
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19107 12804 19717 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20622 12832 20628 12844
rect 20583 12804 20628 12832
rect 20165 12795 20223 12801
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 12124 12736 14841 12764
rect 12124 12724 12130 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 15010 12764 15016 12776
rect 14971 12736 15016 12764
rect 14829 12727 14887 12733
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 17586 12764 17592 12776
rect 15344 12736 17172 12764
rect 17547 12736 17592 12764
rect 15344 12724 15350 12736
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 17037 12699 17095 12705
rect 17037 12696 17049 12699
rect 14792 12668 17049 12696
rect 14792 12656 14798 12668
rect 17037 12665 17049 12668
rect 17083 12665 17095 12699
rect 17037 12659 17095 12665
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13170 12628 13176 12640
rect 12943 12600 13176 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 16761 12631 16819 12637
rect 16761 12597 16773 12631
rect 16807 12628 16819 12631
rect 16942 12628 16948 12640
rect 16807 12600 16948 12628
rect 16807 12597 16819 12600
rect 16761 12591 16819 12597
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 17144 12628 17172 12736
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 19076 12736 19165 12764
rect 19076 12708 19104 12736
rect 19153 12733 19165 12736
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19886 12764 19892 12776
rect 19383 12736 19892 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19886 12724 19892 12736
rect 19944 12724 19950 12776
rect 19058 12656 19064 12708
rect 19116 12656 19122 12708
rect 20180 12628 20208 12795
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 20898 12792 20904 12844
rect 20956 12832 20962 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20956 12804 21097 12832
rect 20956 12792 20962 12804
rect 21085 12801 21097 12804
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 21082 12696 21088 12708
rect 20864 12668 21088 12696
rect 20864 12656 20870 12668
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 17144 12600 20208 12628
rect 20349 12631 20407 12637
rect 20349 12597 20361 12631
rect 20395 12628 20407 12631
rect 21358 12628 21364 12640
rect 20395 12600 21364 12628
rect 20395 12597 20407 12600
rect 20349 12591 20407 12597
rect 21358 12588 21364 12600
rect 21416 12588 21422 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 11977 12427 12035 12433
rect 11977 12424 11989 12427
rect 11940 12396 11989 12424
rect 11940 12384 11946 12396
rect 11977 12393 11989 12396
rect 12023 12393 12035 12427
rect 11977 12387 12035 12393
rect 14829 12427 14887 12433
rect 14829 12393 14841 12427
rect 14875 12424 14887 12427
rect 15010 12424 15016 12436
rect 14875 12396 15016 12424
rect 14875 12393 14887 12396
rect 14829 12387 14887 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15120 12396 15700 12424
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12356 10563 12359
rect 13630 12356 13636 12368
rect 10551 12328 13636 12356
rect 10551 12325 10563 12328
rect 10505 12319 10563 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 15120 12356 15148 12396
rect 13780 12328 15148 12356
rect 15672 12356 15700 12396
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 16264 12396 16313 12424
rect 16264 12384 16270 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 18966 12384 18972 12436
rect 19024 12424 19030 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 19024 12396 19257 12424
rect 19024 12384 19030 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 19702 12384 19708 12436
rect 19760 12424 19766 12436
rect 20625 12427 20683 12433
rect 20625 12424 20637 12427
rect 19760 12396 20637 12424
rect 19760 12384 19766 12396
rect 20625 12393 20637 12396
rect 20671 12393 20683 12427
rect 21266 12424 21272 12436
rect 21227 12396 21272 12424
rect 20625 12387 20683 12393
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 15672 12328 15976 12356
rect 13780 12316 13786 12328
rect 9858 12288 9864 12300
rect 9819 12260 9864 12288
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 11238 12248 11244 12300
rect 11296 12288 11302 12300
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 11296 12260 12541 12288
rect 11296 12248 11302 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 13320 12260 13553 12288
rect 13320 12248 13326 12260
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 13872 12260 14197 12288
rect 13872 12248 13878 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 15838 12288 15844 12300
rect 15799 12260 15844 12288
rect 14185 12251 14243 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 15948 12288 15976 12328
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 17494 12356 17500 12368
rect 17000 12328 17500 12356
rect 17000 12316 17006 12328
rect 17494 12316 17500 12328
rect 17552 12356 17558 12368
rect 18785 12359 18843 12365
rect 18785 12356 18797 12359
rect 17552 12328 18797 12356
rect 17552 12316 17558 12328
rect 18785 12325 18797 12328
rect 18831 12325 18843 12359
rect 18785 12319 18843 12325
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 15948 12260 16865 12288
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17092 12260 17877 12288
rect 17092 12248 17098 12260
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 12437 12223 12495 12229
rect 7892 12192 10916 12220
rect 7892 12180 7898 12192
rect 10137 12155 10195 12161
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 10183 12124 10793 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 10888 12152 10916 12192
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 12483 12192 14381 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 14369 12189 14381 12192
rect 14415 12220 14427 12223
rect 15470 12220 15476 12232
rect 14415 12192 15476 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 16390 12220 16396 12232
rect 15703 12192 16396 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12220 16819 12223
rect 16807 12192 17908 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 10888 12124 13032 12152
rect 10781 12115 10839 12121
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 13004 12093 13032 12124
rect 13814 12112 13820 12164
rect 13872 12152 13878 12164
rect 14461 12155 14519 12161
rect 14461 12152 14473 12155
rect 13872 12124 14473 12152
rect 13872 12112 13878 12124
rect 14461 12121 14473 12124
rect 14507 12121 14519 12155
rect 14461 12115 14519 12121
rect 15749 12155 15807 12161
rect 15749 12121 15761 12155
rect 15795 12152 15807 12155
rect 17880 12152 17908 12192
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 18012 12192 18337 12220
rect 18012 12180 18018 12192
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18800 12220 18828 12319
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 21082 12356 21088 12368
rect 20956 12328 21088 12356
rect 20956 12316 20962 12328
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 20254 12288 20260 12300
rect 19935 12260 20260 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 18800 12192 19625 12220
rect 18325 12183 18383 12189
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19518 12152 19524 12164
rect 15795 12124 17356 12152
rect 17880 12124 19524 12152
rect 15795 12121 15807 12124
rect 15749 12115 15807 12121
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 11296 12056 11621 12084
rect 11296 12044 11302 12056
rect 11609 12053 11621 12056
rect 11655 12084 11667 12087
rect 12345 12087 12403 12093
rect 12345 12084 12357 12087
rect 11655 12056 12357 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 12345 12053 12357 12056
rect 12391 12053 12403 12087
rect 12345 12047 12403 12053
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 13228 12056 13369 12084
rect 13228 12044 13234 12056
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 13357 12047 13415 12053
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 15194 12084 15200 12096
rect 13495 12056 15200 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15289 12087 15347 12093
rect 15289 12053 15301 12087
rect 15335 12084 15347 12087
rect 15378 12084 15384 12096
rect 15335 12056 15384 12084
rect 15335 12053 15347 12056
rect 15289 12047 15347 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 17328 12093 17356 12124
rect 19518 12112 19524 12124
rect 19576 12112 19582 12164
rect 19628 12152 19656 12183
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 20809 12223 20867 12229
rect 20809 12220 20821 12223
rect 20128 12192 20821 12220
rect 20128 12180 20134 12192
rect 20809 12189 20821 12192
rect 20855 12189 20867 12223
rect 21082 12220 21088 12232
rect 21043 12192 21088 12220
rect 20809 12183 20867 12189
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 20257 12155 20315 12161
rect 20257 12152 20269 12155
rect 19628 12124 20269 12152
rect 20257 12121 20269 12124
rect 20303 12121 20315 12155
rect 20257 12115 20315 12121
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 16080 12056 16681 12084
rect 16080 12044 16086 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16669 12047 16727 12053
rect 17313 12087 17371 12093
rect 17313 12053 17325 12087
rect 17359 12053 17371 12087
rect 17313 12047 17371 12053
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 17681 12087 17739 12093
rect 17681 12084 17693 12087
rect 17552 12056 17693 12084
rect 17552 12044 17558 12056
rect 17681 12053 17693 12056
rect 17727 12053 17739 12087
rect 17681 12047 17739 12053
rect 17773 12087 17831 12093
rect 17773 12053 17785 12087
rect 17819 12084 17831 12087
rect 18414 12084 18420 12096
rect 17819 12056 18420 12084
rect 17819 12053 17831 12056
rect 17773 12047 17831 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18509 12087 18567 12093
rect 18509 12053 18521 12087
rect 18555 12084 18567 12087
rect 18598 12084 18604 12096
rect 18555 12056 18604 12084
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 19794 12084 19800 12096
rect 19751 12056 19800 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 9364 11852 11989 11880
rect 9364 11840 9370 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 15286 11880 15292 11892
rect 15247 11852 15292 11880
rect 11977 11843 12035 11849
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 17586 11880 17592 11892
rect 15528 11852 17592 11880
rect 15528 11840 15534 11852
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 17681 11883 17739 11889
rect 17681 11849 17693 11883
rect 17727 11880 17739 11883
rect 18233 11883 18291 11889
rect 18233 11880 18245 11883
rect 17727 11852 18245 11880
rect 17727 11849 17739 11852
rect 17681 11843 17739 11849
rect 18233 11849 18245 11852
rect 18279 11849 18291 11883
rect 18233 11843 18291 11849
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19245 11883 19303 11889
rect 19245 11880 19257 11883
rect 19116 11852 19257 11880
rect 19116 11840 19122 11852
rect 19245 11849 19257 11852
rect 19291 11849 19303 11883
rect 19245 11843 19303 11849
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19702 11880 19708 11892
rect 19576 11852 19708 11880
rect 19576 11840 19582 11852
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11849 20499 11883
rect 20441 11843 20499 11849
rect 21177 11883 21235 11889
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 21450 11880 21456 11892
rect 21223 11852 21456 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 2041 11815 2099 11821
rect 2041 11781 2053 11815
rect 2087 11812 2099 11815
rect 2087 11784 12756 11812
rect 2087 11781 2099 11784
rect 2041 11775 2099 11781
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2056 11744 2084 11775
rect 1719 11716 2084 11744
rect 11701 11747 11759 11753
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 12342 11744 12348 11756
rect 11747 11716 12348 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12618 11676 12624 11688
rect 12492 11648 12537 11676
rect 12579 11648 12624 11676
rect 12492 11636 12498 11648
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 12728 11608 12756 11784
rect 13630 11772 13636 11824
rect 13688 11812 13694 11824
rect 13688 11784 20300 11812
rect 13688 11772 13694 11784
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 14967 11716 15577 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15712 11716 16681 11744
rect 15712 11704 15718 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 18046 11744 18052 11756
rect 17635 11716 18052 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 19610 11744 19616 11756
rect 19571 11716 19616 11744
rect 18601 11707 18659 11713
rect 12802 11636 12808 11688
rect 12860 11676 12866 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 12860 11648 14657 11676
rect 12860 11636 12866 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 14645 11639 14703 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 17736 11648 17785 11676
rect 17736 11636 17742 11648
rect 17773 11645 17785 11648
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 16942 11608 16948 11620
rect 12728 11580 16948 11608
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17494 11568 17500 11620
rect 17552 11608 17558 11620
rect 18616 11608 18644 11707
rect 19610 11704 19616 11716
rect 19668 11704 19674 11756
rect 20272 11753 20300 11784
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11713 20315 11747
rect 20456 11744 20484 11843
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 20772 11784 21404 11812
rect 20772 11772 20778 11784
rect 21376 11753 21404 11784
rect 20901 11747 20959 11753
rect 20901 11744 20913 11747
rect 20456 11716 20913 11744
rect 20257 11707 20315 11713
rect 20901 11713 20913 11716
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 21361 11747 21419 11753
rect 21361 11713 21373 11747
rect 21407 11713 21419 11747
rect 21361 11707 21419 11713
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 17552 11580 18644 11608
rect 18708 11608 18736 11639
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 19889 11679 19947 11685
rect 18840 11648 18885 11676
rect 18840 11636 18846 11648
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 19978 11676 19984 11688
rect 19935 11648 19984 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 21266 11676 21272 11688
rect 20364 11648 21272 11676
rect 20364 11608 20392 11648
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 18708 11580 20392 11608
rect 17552 11568 17558 11580
rect 20438 11568 20444 11620
rect 20496 11608 20502 11620
rect 20717 11611 20775 11617
rect 20717 11608 20729 11611
rect 20496 11580 20729 11608
rect 20496 11568 20502 11580
rect 20717 11577 20729 11580
rect 20763 11577 20775 11611
rect 20717 11571 20775 11577
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16117 11543 16175 11549
rect 16117 11540 16129 11543
rect 16080 11512 16129 11540
rect 16080 11500 16086 11512
rect 16117 11509 16129 11512
rect 16163 11509 16175 11543
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 16117 11503 16175 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 17092 11512 17233 11540
rect 17092 11500 17098 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 22186 11540 22192 11552
rect 19576 11512 22192 11540
rect 19576 11500 19582 11512
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14884 11308 14933 11336
rect 14884 11296 14890 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 14921 11299 14979 11305
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 17678 11336 17684 11348
rect 17359 11308 17684 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 17773 11339 17831 11345
rect 17773 11305 17785 11339
rect 17819 11336 17831 11339
rect 17862 11336 17868 11348
rect 17819 11308 17868 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 18472 11308 18705 11336
rect 18472 11296 18478 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 19518 11336 19524 11348
rect 19479 11308 19524 11336
rect 18693 11299 18751 11305
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 19794 11336 19800 11348
rect 19755 11308 19800 11336
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20257 11339 20315 11345
rect 20257 11336 20269 11339
rect 20036 11308 20269 11336
rect 20036 11296 20042 11308
rect 20257 11305 20269 11308
rect 20303 11305 20315 11339
rect 20257 11299 20315 11305
rect 20717 11339 20775 11345
rect 20717 11305 20729 11339
rect 20763 11336 20775 11339
rect 21174 11336 21180 11348
rect 20763 11308 21036 11336
rect 21135 11308 21180 11336
rect 20763 11305 20775 11308
rect 20717 11299 20775 11305
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 12492 11240 14504 11268
rect 12492 11228 12498 11240
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 14476 11209 14504 11240
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 21008 11268 21036 11308
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 21634 11268 21640 11280
rect 16908 11240 20944 11268
rect 21008 11240 21640 11268
rect 16908 11228 16914 11240
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 11756 11172 14289 11200
rect 11756 11160 11762 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 15838 11200 15844 11212
rect 14507 11172 15844 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16025 11203 16083 11209
rect 16025 11169 16037 11203
rect 16071 11200 16083 11203
rect 18046 11200 18052 11212
rect 16071 11172 17908 11200
rect 18007 11172 18052 11200
rect 16071 11169 16083 11172
rect 16025 11163 16083 11169
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11101 17187 11135
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17129 11095 17187 11101
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 14553 11067 14611 11073
rect 14553 11064 14565 11067
rect 7340 11036 14565 11064
rect 7340 11024 7346 11036
rect 14553 11033 14565 11036
rect 14599 11033 14611 11067
rect 14553 11027 14611 11033
rect 16393 11067 16451 11073
rect 16393 11033 16405 11067
rect 16439 11064 16451 11067
rect 17144 11064 17172 11095
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 17880 11132 17908 11172
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 19058 11200 19064 11212
rect 18800 11172 19064 11200
rect 18800 11132 18828 11172
rect 19058 11160 19064 11172
rect 19116 11200 19122 11212
rect 19116 11172 20484 11200
rect 19116 11160 19122 11172
rect 17880 11104 18828 11132
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 19334 11132 19340 11144
rect 19295 11104 19340 11132
rect 18877 11095 18935 11101
rect 17954 11064 17960 11076
rect 16439 11036 17960 11064
rect 16439 11033 16451 11036
rect 16393 11027 16451 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 18892 11064 18920 11095
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19978 11132 19984 11144
rect 19891 11104 19984 11132
rect 19978 11092 19984 11104
rect 20036 11132 20042 11144
rect 20254 11132 20260 11144
rect 20036 11104 20260 11132
rect 20036 11092 20042 11104
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 20456 11141 20484 11172
rect 20916 11141 20944 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11101 20499 11135
rect 20441 11095 20499 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 21358 11132 21364 11144
rect 21319 11104 21364 11132
rect 20901 11095 20959 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 21450 11064 21456 11076
rect 18892 11036 21456 11064
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 15286 10996 15292 11008
rect 15247 10968 15292 10996
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 16669 10999 16727 11005
rect 16669 10965 16681 10999
rect 16715 10996 16727 10999
rect 16942 10996 16948 11008
rect 16715 10968 16948 10996
rect 16715 10965 16727 10968
rect 16669 10959 16727 10965
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15286 10792 15292 10804
rect 15243 10764 15292 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15565 10795 15623 10801
rect 15565 10761 15577 10795
rect 15611 10792 15623 10795
rect 15654 10792 15660 10804
rect 15611 10764 15660 10792
rect 15611 10761 15623 10764
rect 15565 10755 15623 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 17310 10752 17316 10804
rect 17368 10752 17374 10804
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10761 17739 10795
rect 17681 10755 17739 10761
rect 18141 10795 18199 10801
rect 18141 10761 18153 10795
rect 18187 10792 18199 10795
rect 18506 10792 18512 10804
rect 18187 10764 18512 10792
rect 18187 10761 18199 10764
rect 18141 10755 18199 10761
rect 17328 10724 17356 10752
rect 14936 10696 17356 10724
rect 14936 10597 14964 10696
rect 17310 10656 17316 10668
rect 17271 10628 17316 10656
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17696 10656 17724 10755
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 18601 10795 18659 10801
rect 18601 10761 18613 10795
rect 18647 10792 18659 10795
rect 19334 10792 19340 10804
rect 18647 10764 19340 10792
rect 18647 10761 18659 10764
rect 18601 10755 18659 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10761 20131 10795
rect 20530 10792 20536 10804
rect 20491 10764 20536 10792
rect 20073 10755 20131 10761
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 20088 10724 20116 10755
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 20806 10752 20812 10804
rect 20864 10752 20870 10804
rect 20990 10792 20996 10804
rect 20951 10764 20996 10792
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 21361 10795 21419 10801
rect 21361 10761 21373 10795
rect 21407 10792 21419 10795
rect 21450 10792 21456 10804
rect 21407 10764 21456 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 20824 10724 20852 10752
rect 17920 10696 18920 10724
rect 20088 10696 20852 10724
rect 17920 10684 17926 10696
rect 17957 10659 18015 10665
rect 17957 10656 17969 10659
rect 17696 10628 17969 10656
rect 17957 10625 17969 10628
rect 18003 10625 18015 10659
rect 17957 10619 18015 10625
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 18690 10656 18696 10668
rect 18463 10628 18696 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 18892 10665 18920 10696
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 19429 10659 19487 10665
rect 19429 10625 19441 10659
rect 19475 10625 19487 10659
rect 19886 10656 19892 10668
rect 19847 10628 19892 10656
rect 19429 10619 19487 10625
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 15068 10560 15117 10588
rect 15068 10548 15074 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 17126 10588 17132 10600
rect 17087 10560 17132 10588
rect 15105 10551 15163 10557
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10557 17279 10591
rect 17221 10551 17279 10557
rect 17236 10520 17264 10551
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 19444 10588 19472 10619
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 20346 10656 20352 10668
rect 20307 10628 20352 10656
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 18656 10560 19472 10588
rect 18656 10548 18662 10560
rect 17954 10520 17960 10532
rect 17236 10492 17960 10520
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 19061 10523 19119 10529
rect 19061 10489 19073 10523
rect 19107 10520 19119 10523
rect 20622 10520 20628 10532
rect 19107 10492 20628 10520
rect 19107 10489 19119 10492
rect 19061 10483 19119 10489
rect 20622 10480 20628 10492
rect 20680 10480 20686 10532
rect 15930 10412 15936 10464
rect 15988 10452 15994 10464
rect 19518 10452 19524 10464
rect 15988 10424 19524 10452
rect 15988 10412 15994 10424
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19613 10455 19671 10461
rect 19613 10421 19625 10455
rect 19659 10452 19671 10455
rect 22370 10452 22376 10464
rect 19659 10424 22376 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 17037 10251 17095 10257
rect 17037 10217 17049 10251
rect 17083 10248 17095 10251
rect 17586 10248 17592 10260
rect 17083 10220 17592 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18690 10248 18696 10260
rect 18651 10220 18696 10248
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19613 10251 19671 10257
rect 19613 10217 19625 10251
rect 19659 10248 19671 10251
rect 20806 10248 20812 10260
rect 19659 10220 20812 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 15930 10180 15936 10192
rect 11204 10152 15936 10180
rect 11204 10140 11210 10152
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 20070 10180 20076 10192
rect 17276 10152 18092 10180
rect 20031 10152 20076 10180
rect 17276 10140 17282 10152
rect 15562 10112 15568 10124
rect 15523 10084 15568 10112
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10112 16543 10115
rect 17402 10112 17408 10124
rect 16531 10084 17408 10112
rect 16531 10081 16543 10084
rect 16485 10075 16543 10081
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 18064 10121 18092 10152
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 20349 10183 20407 10189
rect 20349 10149 20361 10183
rect 20395 10149 20407 10183
rect 20349 10143 20407 10149
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15470 10044 15476 10056
rect 15252 10016 15476 10044
rect 15252 10004 15258 10016
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10044 16727 10047
rect 16942 10044 16948 10056
rect 16715 10016 16948 10044
rect 16715 10013 16727 10016
rect 16669 10007 16727 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17494 10004 17500 10056
rect 17552 10044 17558 10056
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 17552 10016 17693 10044
rect 17552 10004 17558 10016
rect 17681 10013 17693 10016
rect 17727 10044 17739 10047
rect 18230 10044 18236 10056
rect 17727 10016 18236 10044
rect 17727 10013 17739 10016
rect 17681 10007 17739 10013
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20364 10044 20392 10143
rect 20993 10115 21051 10121
rect 20993 10081 21005 10115
rect 21039 10112 21051 10115
rect 22738 10112 22744 10124
rect 21039 10084 22744 10112
rect 21039 10081 21051 10084
rect 20993 10075 21051 10081
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 19935 10016 20392 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 8168 9948 15393 9976
rect 8168 9936 8174 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15381 9939 15439 9945
rect 16577 9979 16635 9985
rect 16577 9945 16589 9979
rect 16623 9976 16635 9979
rect 17218 9976 17224 9988
rect 16623 9948 17224 9976
rect 16623 9945 16635 9948
rect 16577 9939 16635 9945
rect 17218 9936 17224 9948
rect 17276 9936 17282 9988
rect 19444 9976 19472 10007
rect 20162 9976 20168 9988
rect 19444 9948 20168 9976
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 14737 9911 14795 9917
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 15194 9908 15200 9920
rect 14783 9880 15200 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 15194 9868 15200 9880
rect 15252 9868 15258 9920
rect 16942 9868 16948 9920
rect 17000 9908 17006 9920
rect 17497 9911 17555 9917
rect 17497 9908 17509 9911
rect 17000 9880 17509 9908
rect 17000 9868 17006 9880
rect 17497 9877 17509 9880
rect 17543 9877 17555 9911
rect 18230 9908 18236 9920
rect 18191 9880 18236 9908
rect 17497 9871 17555 9877
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18322 9868 18328 9920
rect 18380 9908 18386 9920
rect 20714 9908 20720 9920
rect 18380 9880 18425 9908
rect 20675 9880 20720 9908
rect 18380 9868 18386 9880
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20809 9911 20867 9917
rect 20809 9877 20821 9911
rect 20855 9908 20867 9911
rect 20990 9908 20996 9920
rect 20855 9880 20996 9908
rect 20855 9877 20867 9880
rect 20809 9871 20867 9877
rect 20990 9868 20996 9880
rect 21048 9868 21054 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 17494 9704 17500 9716
rect 17455 9676 17500 9704
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 18230 9704 18236 9716
rect 18191 9676 18236 9704
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18693 9707 18751 9713
rect 18693 9673 18705 9707
rect 18739 9704 18751 9707
rect 19705 9707 19763 9713
rect 18739 9676 18920 9704
rect 18739 9673 18751 9676
rect 18693 9667 18751 9673
rect 11790 9596 11796 9648
rect 11848 9636 11854 9648
rect 15194 9636 15200 9648
rect 11848 9608 12756 9636
rect 15155 9608 15200 9636
rect 11848 9596 11854 9608
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12728 9509 12756 9608
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 18892 9636 18920 9676
rect 19705 9673 19717 9707
rect 19751 9704 19763 9707
rect 19886 9704 19892 9716
rect 19751 9676 19892 9704
rect 19751 9673 19763 9676
rect 19705 9667 19763 9673
rect 19886 9664 19892 9676
rect 19944 9664 19950 9716
rect 20162 9704 20168 9716
rect 20123 9676 20168 9704
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 19610 9636 19616 9648
rect 18892 9608 19616 9636
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 17770 9568 17776 9580
rect 17731 9540 17776 9568
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18230 9528 18236 9580
rect 18288 9568 18294 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18288 9540 18613 9568
rect 18288 9528 18294 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 19518 9568 19524 9580
rect 19479 9540 19524 9568
rect 18601 9531 18659 9537
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9568 21419 9571
rect 21634 9568 21640 9580
rect 21407 9540 21640 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9469 12771 9503
rect 12713 9463 12771 9469
rect 12158 9432 12164 9444
rect 12119 9404 12164 9432
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12636 9432 12664 9463
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 12952 9472 14933 9500
rect 12952 9460 12958 9472
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 15105 9503 15163 9509
rect 15105 9469 15117 9503
rect 15151 9500 15163 9503
rect 15562 9500 15568 9512
rect 15151 9472 15568 9500
rect 15151 9469 15163 9472
rect 15105 9463 15163 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 18414 9460 18420 9512
rect 18472 9500 18478 9512
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 18472 9472 18797 9500
rect 18472 9460 18478 9472
rect 18785 9469 18797 9472
rect 18831 9469 18843 9503
rect 20622 9500 20628 9512
rect 20583 9472 20628 9500
rect 18785 9463 18843 9469
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9500 20867 9503
rect 20898 9500 20904 9512
rect 20855 9472 20904 9500
rect 20855 9469 20867 9472
rect 20809 9463 20867 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 15010 9432 15016 9444
rect 12636 9404 15016 9432
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 17862 9432 17868 9444
rect 15580 9404 17868 9432
rect 15580 9373 15608 9404
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 17957 9435 18015 9441
rect 17957 9401 17969 9435
rect 18003 9432 18015 9435
rect 20346 9432 20352 9444
rect 18003 9404 20352 9432
rect 18003 9401 18015 9404
rect 17957 9395 18015 9401
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 21376 9432 21404 9531
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 20456 9404 21404 9432
rect 15565 9367 15623 9373
rect 15565 9333 15577 9367
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 20456 9364 20484 9404
rect 21174 9364 21180 9376
rect 17175 9336 20484 9364
rect 21135 9336 21180 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 15562 9160 15568 9172
rect 15523 9132 15568 9160
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9160 17003 9163
rect 17310 9160 17316 9172
rect 16991 9132 17316 9160
rect 16991 9129 17003 9132
rect 16945 9123 17003 9129
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17957 9163 18015 9169
rect 17957 9129 17969 9163
rect 18003 9160 18015 9163
rect 18322 9160 18328 9172
rect 18003 9132 18328 9160
rect 18003 9129 18015 9132
rect 17957 9123 18015 9129
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 19337 9163 19395 9169
rect 19337 9129 19349 9163
rect 19383 9160 19395 9163
rect 19978 9160 19984 9172
rect 19383 9132 19984 9160
rect 19383 9129 19395 9132
rect 19337 9123 19395 9129
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20622 9120 20628 9172
rect 20680 9160 20686 9172
rect 20809 9163 20867 9169
rect 20809 9160 20821 9163
rect 20680 9132 20821 9160
rect 20680 9120 20686 9132
rect 20809 9129 20821 9132
rect 20855 9129 20867 9163
rect 21082 9160 21088 9172
rect 21043 9132 21088 9160
rect 20809 9123 20867 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 15838 9052 15844 9104
rect 15896 9092 15902 9104
rect 19797 9095 19855 9101
rect 15896 9064 19564 9092
rect 15896 9052 15902 9064
rect 15013 9027 15071 9033
rect 15013 8993 15025 9027
rect 15059 9024 15071 9027
rect 16114 9024 16120 9036
rect 15059 8996 16120 9024
rect 15059 8993 15071 8996
rect 15013 8987 15071 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16298 9024 16304 9036
rect 16259 8996 16304 9024
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 18414 9024 18420 9036
rect 17451 8996 18420 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 12406 8928 15853 8956
rect 12406 8888 12434 8928
rect 15841 8925 15853 8928
rect 15887 8956 15899 8959
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 15887 8928 16497 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 18322 8956 18328 8968
rect 16485 8919 16543 8925
rect 17512 8928 18328 8956
rect 15197 8891 15255 8897
rect 15197 8888 15209 8891
rect 6886 8860 12434 8888
rect 13464 8860 15209 8888
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 6886 8820 6914 8860
rect 5132 8792 6914 8820
rect 5132 8780 5138 8792
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 13464 8820 13492 8860
rect 15197 8857 15209 8860
rect 15243 8857 15255 8891
rect 17512 8888 17540 8928
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8956 18935 8959
rect 18966 8956 18972 8968
rect 18923 8928 18972 8956
rect 18923 8925 18935 8928
rect 18877 8919 18935 8925
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 15197 8851 15255 8857
rect 16500 8860 17540 8888
rect 17589 8891 17647 8897
rect 7708 8792 13492 8820
rect 7708 8780 7714 8792
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15105 8823 15163 8829
rect 15105 8820 15117 8823
rect 15068 8792 15117 8820
rect 15068 8780 15074 8792
rect 15105 8789 15117 8792
rect 15151 8820 15163 8823
rect 16500 8820 16528 8860
rect 17589 8857 17601 8891
rect 17635 8888 17647 8891
rect 18233 8891 18291 8897
rect 18233 8888 18245 8891
rect 17635 8860 18245 8888
rect 17635 8857 17647 8860
rect 17589 8851 17647 8857
rect 18233 8857 18245 8860
rect 18279 8857 18291 8891
rect 19536 8888 19564 9064
rect 19797 9061 19809 9095
rect 19843 9061 19855 9095
rect 19797 9055 19855 9061
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8956 19671 8959
rect 19702 8956 19708 8968
rect 19659 8928 19708 8956
rect 19659 8925 19671 8928
rect 19613 8919 19671 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 19812 8956 19840 9055
rect 19886 8984 19892 9036
rect 19944 9024 19950 9036
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 19944 8996 20177 9024
rect 19944 8984 19950 8996
rect 20165 8993 20177 8996
rect 20211 9024 20223 9027
rect 20898 9024 20904 9036
rect 20211 8996 20904 9024
rect 20211 8993 20223 8996
rect 20165 8987 20223 8993
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 19812 8928 21281 8956
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 20622 8888 20628 8900
rect 19536 8860 20628 8888
rect 18233 8851 18291 8857
rect 20622 8848 20628 8860
rect 20680 8848 20686 8900
rect 15151 8792 16528 8820
rect 16577 8823 16635 8829
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 16577 8789 16589 8823
rect 16623 8820 16635 8823
rect 17126 8820 17132 8832
rect 16623 8792 17132 8820
rect 16623 8789 16635 8792
rect 16577 8783 16635 8789
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 17494 8820 17500 8832
rect 17455 8792 17500 8820
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18693 8823 18751 8829
rect 18693 8820 18705 8823
rect 18104 8792 18705 8820
rect 18104 8780 18110 8792
rect 18693 8789 18705 8792
rect 18739 8789 18751 8823
rect 18693 8783 18751 8789
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19610 8820 19616 8832
rect 19392 8792 19616 8820
rect 19392 8780 19398 8792
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 20346 8820 20352 8832
rect 20307 8792 20352 8820
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20441 8823 20499 8829
rect 20441 8789 20453 8823
rect 20487 8820 20499 8823
rect 20806 8820 20812 8832
rect 20487 8792 20812 8820
rect 20487 8789 20499 8792
rect 20441 8783 20499 8789
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 17954 8616 17960 8628
rect 16347 8588 17816 8616
rect 17915 8588 17960 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 17494 8548 17500 8560
rect 9272 8520 17500 8548
rect 9272 8508 9278 8520
rect 17494 8508 17500 8520
rect 17552 8508 17558 8560
rect 17788 8548 17816 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18417 8619 18475 8625
rect 18417 8585 18429 8619
rect 18463 8616 18475 8619
rect 19334 8616 19340 8628
rect 18463 8588 19340 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19702 8616 19708 8628
rect 19663 8588 19708 8616
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20714 8616 20720 8628
rect 20675 8588 20720 8616
rect 20714 8576 20720 8588
rect 20772 8576 20778 8628
rect 21177 8619 21235 8625
rect 21177 8585 21189 8619
rect 21223 8616 21235 8619
rect 21266 8616 21272 8628
rect 21223 8588 21272 8616
rect 21223 8585 21235 8588
rect 21177 8579 21235 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 20073 8551 20131 8557
rect 17788 8520 20024 8548
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 17126 8480 17132 8492
rect 16715 8452 17132 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17267 8452 17693 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17681 8449 17693 8452
rect 17727 8480 17739 8483
rect 17954 8480 17960 8492
rect 17727 8452 17960 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 18288 8452 18337 8480
rect 18288 8440 18294 8452
rect 18325 8449 18337 8452
rect 18371 8480 18383 8483
rect 18371 8452 18644 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 16298 8372 16304 8424
rect 16356 8412 16362 8424
rect 18509 8415 18567 8421
rect 16356 8384 18368 8412
rect 16356 8372 16362 8384
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 16172 8316 17509 8344
rect 16172 8304 16178 8316
rect 17497 8313 17509 8316
rect 17543 8313 17555 8347
rect 18340 8344 18368 8384
rect 18509 8381 18521 8415
rect 18555 8381 18567 8415
rect 18616 8412 18644 8452
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 19242 8480 19248 8492
rect 18840 8452 19248 8480
rect 18840 8440 18846 8452
rect 19242 8440 19248 8452
rect 19300 8480 19306 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19300 8452 19441 8480
rect 19300 8440 19306 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19996 8480 20024 8520
rect 20073 8517 20085 8551
rect 20119 8548 20131 8551
rect 20254 8548 20260 8560
rect 20119 8520 20260 8548
rect 20119 8517 20131 8520
rect 20073 8511 20131 8517
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 21358 8480 21364 8492
rect 19996 8452 21364 8480
rect 19429 8443 19487 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 20162 8412 20168 8424
rect 18616 8384 19380 8412
rect 20123 8384 20168 8412
rect 18509 8375 18567 8381
rect 18524 8344 18552 8375
rect 18340 8316 18552 8344
rect 17497 8307 17555 8313
rect 18690 8304 18696 8356
rect 18748 8344 18754 8356
rect 19245 8347 19303 8353
rect 19245 8344 19257 8347
rect 18748 8316 19257 8344
rect 18748 8304 18754 8316
rect 19245 8313 19257 8316
rect 19291 8313 19303 8347
rect 19352 8344 19380 8384
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8412 20407 8415
rect 22094 8412 22100 8424
rect 20395 8384 22100 8412
rect 20395 8381 20407 8384
rect 20349 8375 20407 8381
rect 22094 8372 22100 8384
rect 22152 8372 22158 8424
rect 21266 8344 21272 8356
rect 19352 8316 21272 8344
rect 19245 8307 19303 8313
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 19886 8276 19892 8288
rect 15528 8248 19892 8276
rect 15528 8236 15534 8248
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 17770 8072 17776 8084
rect 17727 8044 17776 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18782 8072 18788 8084
rect 18616 8044 18788 8072
rect 17037 8007 17095 8013
rect 17037 7973 17049 8007
rect 17083 8004 17095 8007
rect 18616 8004 18644 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 20346 8072 20352 8084
rect 20307 8044 20352 8072
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 17083 7976 18644 8004
rect 17083 7973 17095 7976
rect 17037 7967 17095 7973
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 21174 8004 21180 8016
rect 18748 7976 21180 8004
rect 18748 7964 18754 7976
rect 21174 7964 21180 7976
rect 21232 7964 21238 8016
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 18233 7939 18291 7945
rect 18233 7936 18245 7939
rect 18196 7908 18245 7936
rect 18196 7896 18202 7908
rect 18233 7905 18245 7908
rect 18279 7905 18291 7939
rect 18233 7899 18291 7905
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 19610 7936 19616 7948
rect 19567 7908 19616 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 19610 7896 19616 7908
rect 19668 7936 19674 7948
rect 20070 7936 20076 7948
rect 19668 7908 20076 7936
rect 19668 7896 19674 7908
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20772 7908 21005 7936
rect 20772 7896 20778 7908
rect 20993 7905 21005 7908
rect 21039 7936 21051 7939
rect 22278 7936 22284 7948
rect 21039 7908 22284 7936
rect 21039 7905 21051 7908
rect 20993 7899 21051 7905
rect 22278 7896 22284 7908
rect 22336 7896 22342 7948
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7868 17463 7871
rect 18877 7871 18935 7877
rect 18877 7868 18889 7871
rect 17451 7840 18889 7868
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 18877 7837 18889 7840
rect 18923 7868 18935 7871
rect 18966 7868 18972 7880
rect 18923 7840 18972 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19702 7868 19708 7880
rect 19615 7840 19708 7868
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 19628 7809 19656 7840
rect 19702 7828 19708 7840
rect 19760 7868 19766 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 19760 7840 20821 7868
rect 19760 7828 19766 7840
rect 20809 7837 20821 7840
rect 20855 7868 20867 7871
rect 22462 7868 22468 7880
rect 20855 7840 22468 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 22462 7828 22468 7840
rect 22520 7828 22526 7880
rect 18049 7803 18107 7809
rect 18049 7800 18061 7803
rect 16356 7772 18061 7800
rect 16356 7760 16362 7772
rect 18049 7769 18061 7772
rect 18095 7769 18107 7803
rect 18049 7763 18107 7769
rect 19613 7803 19671 7809
rect 19613 7769 19625 7803
rect 19659 7769 19671 7803
rect 20717 7803 20775 7809
rect 20717 7800 20729 7803
rect 19613 7763 19671 7769
rect 19904 7772 20729 7800
rect 19904 7744 19932 7772
rect 20717 7769 20729 7772
rect 20763 7769 20775 7803
rect 20717 7763 20775 7769
rect 18138 7692 18144 7744
rect 18196 7732 18202 7744
rect 18196 7704 18241 7732
rect 18196 7692 18202 7704
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 18472 7704 18705 7732
rect 18472 7692 18478 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 18693 7695 18751 7701
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 19886 7732 19892 7744
rect 19751 7704 19892 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 20070 7732 20076 7744
rect 20031 7704 20076 7732
rect 20070 7692 20076 7704
rect 20128 7692 20134 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 15804 7500 17049 7528
rect 15804 7488 15810 7500
rect 17037 7497 17049 7500
rect 17083 7528 17095 7531
rect 17862 7528 17868 7540
rect 17083 7500 17868 7528
rect 17083 7497 17095 7500
rect 17037 7491 17095 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 19337 7531 19395 7537
rect 19337 7497 19349 7531
rect 19383 7528 19395 7531
rect 19518 7528 19524 7540
rect 19383 7500 19524 7528
rect 19383 7497 19395 7500
rect 19337 7491 19395 7497
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 19702 7488 19708 7540
rect 19760 7528 19766 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 19760 7500 20361 7528
rect 19760 7488 19766 7500
rect 20349 7497 20361 7500
rect 20395 7497 20407 7531
rect 20349 7491 20407 7497
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 20806 7528 20812 7540
rect 20763 7500 20812 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 15286 7420 15292 7472
rect 15344 7460 15350 7472
rect 18414 7460 18420 7472
rect 15344 7432 18420 7460
rect 15344 7420 15350 7432
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 18874 7460 18880 7472
rect 18708 7432 18880 7460
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 18322 7392 18328 7404
rect 17911 7364 18328 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 15562 7284 15568 7336
rect 15620 7324 15626 7336
rect 18046 7324 18052 7336
rect 15620 7296 18052 7324
rect 15620 7284 15626 7296
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18708 7333 18736 7432
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 19058 7420 19064 7472
rect 19116 7460 19122 7472
rect 19613 7463 19671 7469
rect 19613 7460 19625 7463
rect 19116 7432 19625 7460
rect 19116 7420 19122 7432
rect 19613 7429 19625 7432
rect 19659 7429 19671 7463
rect 19613 7423 19671 7429
rect 20088 7432 21404 7460
rect 18782 7352 18788 7404
rect 18840 7392 18846 7404
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18840 7364 18981 7392
rect 18840 7352 18846 7364
rect 18969 7361 18981 7364
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18874 7324 18880 7336
rect 18835 7296 18880 7324
rect 18693 7287 18751 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 16761 7259 16819 7265
rect 16761 7225 16773 7259
rect 16807 7256 16819 7259
rect 20088 7256 20116 7432
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20622 7392 20628 7404
rect 20303 7364 20628 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 21376 7401 21404 7432
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21450 7392 21456 7404
rect 21407 7364 21456 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 20165 7327 20223 7333
rect 20165 7293 20177 7327
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 16807 7228 20116 7256
rect 20180 7256 20208 7287
rect 20714 7256 20720 7268
rect 20180 7228 20720 7256
rect 16807 7225 16819 7228
rect 16761 7219 16819 7225
rect 20714 7216 20720 7228
rect 20772 7216 20778 7268
rect 17494 7188 17500 7200
rect 17455 7160 17500 7188
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 18141 7191 18199 7197
rect 18141 7188 18153 7191
rect 18104 7160 18153 7188
rect 18104 7148 18110 7160
rect 18141 7157 18153 7160
rect 18187 7157 18199 7191
rect 21174 7188 21180 7200
rect 21135 7160 21180 7188
rect 18141 7151 18199 7157
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19886 6984 19892 6996
rect 19484 6956 19892 6984
rect 19484 6944 19490 6956
rect 19886 6944 19892 6956
rect 19944 6944 19950 6996
rect 18598 6916 18604 6928
rect 18248 6888 18604 6916
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6848 16911 6851
rect 17310 6848 17316 6860
rect 16899 6820 17316 6848
rect 16899 6817 16911 6820
rect 16853 6811 16911 6817
rect 17052 6712 17080 6820
rect 17310 6808 17316 6820
rect 17368 6848 17374 6860
rect 17586 6848 17592 6860
rect 17368 6820 17592 6848
rect 17368 6808 17374 6820
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 18046 6848 18052 6860
rect 18007 6820 18052 6848
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18248 6857 18276 6888
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 19978 6876 19984 6928
rect 20036 6916 20042 6928
rect 20622 6916 20628 6928
rect 20036 6888 20628 6916
rect 20036 6876 20042 6888
rect 20622 6876 20628 6888
rect 20680 6876 20686 6928
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 19794 6848 19800 6860
rect 19576 6820 19800 6848
rect 19576 6808 19582 6820
rect 19794 6808 19800 6820
rect 19852 6808 19858 6860
rect 19889 6851 19947 6857
rect 19889 6817 19901 6851
rect 19935 6817 19947 6851
rect 19889 6811 19947 6817
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6780 17187 6783
rect 17494 6780 17500 6792
rect 17175 6752 17500 6780
rect 17175 6749 17187 6752
rect 17129 6743 17187 6749
rect 17494 6740 17500 6752
rect 17552 6780 17558 6792
rect 18322 6780 18328 6792
rect 17552 6752 18328 6780
rect 17552 6740 17558 6752
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 18966 6780 18972 6792
rect 18739 6752 18972 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19076 6752 19717 6780
rect 17957 6715 18015 6721
rect 17957 6712 17969 6715
rect 17052 6684 17969 6712
rect 17957 6681 17969 6684
rect 18003 6681 18015 6715
rect 19076 6712 19104 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 17957 6675 18015 6681
rect 18064 6684 19104 6712
rect 17313 6647 17371 6653
rect 17313 6613 17325 6647
rect 17359 6644 17371 6647
rect 17402 6644 17408 6656
rect 17359 6616 17408 6644
rect 17359 6613 17371 6616
rect 17313 6607 17371 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17586 6644 17592 6656
rect 17547 6616 17592 6644
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 18064 6644 18092 6684
rect 19518 6672 19524 6724
rect 19576 6712 19582 6724
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 19576 6684 19625 6712
rect 19576 6672 19582 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 17828 6616 18092 6644
rect 18877 6647 18935 6653
rect 17828 6604 17834 6616
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 18966 6644 18972 6656
rect 18923 6616 18972 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 19242 6644 19248 6656
rect 19203 6616 19248 6644
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19720 6644 19748 6743
rect 19904 6724 19932 6811
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 20128 6820 20729 6848
rect 20128 6808 20134 6820
rect 20717 6817 20729 6820
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 21082 6848 21088 6860
rect 20947 6820 21088 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 21082 6808 21088 6820
rect 21140 6848 21146 6860
rect 21542 6848 21548 6860
rect 21140 6820 21548 6848
rect 21140 6808 21146 6820
rect 21542 6808 21548 6820
rect 21600 6808 21606 6860
rect 19886 6712 19892 6724
rect 19799 6684 19892 6712
rect 19886 6672 19892 6684
rect 19944 6712 19950 6724
rect 21358 6712 21364 6724
rect 19944 6684 20760 6712
rect 21319 6684 21364 6712
rect 19944 6672 19950 6684
rect 20070 6644 20076 6656
rect 19720 6616 20076 6644
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 20162 6604 20168 6656
rect 20220 6644 20226 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 20220 6616 20269 6644
rect 20220 6604 20226 6616
rect 20257 6613 20269 6616
rect 20303 6613 20315 6647
rect 20622 6644 20628 6656
rect 20583 6616 20628 6644
rect 20257 6607 20315 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 20732 6644 20760 6684
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 22646 6644 22652 6656
rect 20732 6616 22652 6644
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 18138 6440 18144 6452
rect 18099 6412 18144 6440
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 19242 6440 19248 6452
rect 18555 6412 19248 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 20349 6443 20407 6449
rect 20349 6409 20361 6443
rect 20395 6440 20407 6443
rect 20530 6440 20536 6452
rect 20395 6412 20536 6440
rect 20395 6409 20407 6412
rect 20349 6403 20407 6409
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 18046 6372 18052 6384
rect 17420 6344 18052 6372
rect 17420 6313 17448 6344
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 19613 6375 19671 6381
rect 19613 6341 19625 6375
rect 19659 6372 19671 6375
rect 20717 6375 20775 6381
rect 20717 6372 20729 6375
rect 19659 6344 20729 6372
rect 19659 6341 19671 6344
rect 19613 6335 19671 6341
rect 20717 6341 20729 6344
rect 20763 6341 20775 6375
rect 20717 6335 20775 6341
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6304 17003 6307
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 16991 6276 17417 6304
rect 16991 6273 17003 6276
rect 16945 6267 17003 6273
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 17770 6304 17776 6316
rect 17552 6276 17776 6304
rect 17552 6264 17558 6276
rect 17770 6264 17776 6276
rect 17828 6264 17834 6316
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 17954 6304 17960 6316
rect 17911 6276 17960 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 17880 6236 17908 6267
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 20073 6307 20131 6313
rect 18564 6276 18736 6304
rect 18564 6264 18570 6276
rect 18598 6236 18604 6248
rect 16347 6208 17908 6236
rect 18559 6208 18604 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 18708 6245 18736 6276
rect 20073 6273 20085 6307
rect 20119 6304 20131 6307
rect 20346 6304 20352 6316
rect 20119 6276 20352 6304
rect 20119 6273 20131 6276
rect 20073 6267 20131 6273
rect 20346 6264 20352 6276
rect 20404 6264 20410 6316
rect 18693 6239 18751 6245
rect 18693 6205 18705 6239
rect 18739 6205 18751 6239
rect 18693 6199 18751 6205
rect 20438 6196 20444 6248
rect 20496 6236 20502 6248
rect 20809 6239 20867 6245
rect 20809 6236 20821 6239
rect 20496 6208 20821 6236
rect 20496 6196 20502 6208
rect 20809 6205 20821 6208
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 20956 6208 21001 6236
rect 20956 6196 20962 6208
rect 10686 6128 10692 6180
rect 10744 6168 10750 6180
rect 13170 6168 13176 6180
rect 10744 6140 13176 6168
rect 10744 6128 10750 6140
rect 13170 6128 13176 6140
rect 13228 6128 13234 6180
rect 15654 6128 15660 6180
rect 15712 6168 15718 6180
rect 17681 6171 17739 6177
rect 17681 6168 17693 6171
rect 15712 6140 17693 6168
rect 15712 6128 15718 6140
rect 17681 6137 17693 6140
rect 17727 6137 17739 6171
rect 17681 6131 17739 6137
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 17221 6103 17279 6109
rect 17221 6100 17233 6103
rect 14884 6072 17233 6100
rect 14884 6060 14890 6072
rect 17221 6069 17233 6072
rect 17267 6069 17279 6103
rect 17221 6063 17279 6069
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 19889 6103 19947 6109
rect 19889 6100 19901 6103
rect 17828 6072 19901 6100
rect 17828 6060 17834 6072
rect 19889 6069 19901 6072
rect 19935 6069 19947 6103
rect 19889 6063 19947 6069
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 14700 5868 17601 5896
rect 14700 5856 14706 5868
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 17589 5859 17647 5865
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 18656 5868 19257 5896
rect 18656 5856 18662 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 20438 5896 20444 5908
rect 20399 5868 20444 5896
rect 19245 5859 19303 5865
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 14366 5788 14372 5840
rect 14424 5828 14430 5840
rect 17129 5831 17187 5837
rect 17129 5828 17141 5831
rect 14424 5800 17141 5828
rect 14424 5788 14430 5800
rect 17129 5797 17141 5800
rect 17175 5797 17187 5831
rect 17862 5828 17868 5840
rect 17129 5791 17187 5797
rect 17236 5800 17868 5828
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 15746 5760 15752 5772
rect 15703 5732 15752 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16439 5664 16865 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16853 5661 16865 5664
rect 16899 5692 16911 5695
rect 17236 5692 17264 5800
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 19886 5760 19892 5772
rect 17460 5732 18460 5760
rect 19847 5732 19892 5760
rect 17460 5720 17466 5732
rect 16899 5664 17264 5692
rect 17313 5695 17371 5701
rect 16899 5661 16911 5664
rect 16853 5655 16911 5661
rect 17313 5661 17325 5695
rect 17359 5661 17371 5695
rect 17313 5655 17371 5661
rect 14274 5584 14280 5636
rect 14332 5624 14338 5636
rect 16025 5627 16083 5633
rect 14332 5596 15700 5624
rect 14332 5584 14338 5596
rect 15672 5556 15700 5596
rect 16025 5593 16037 5627
rect 16071 5624 16083 5627
rect 17328 5624 17356 5655
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17736 5664 17785 5692
rect 17736 5652 17742 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 18432 5701 18460 5732
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20772 5732 21005 5760
rect 20772 5720 20778 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5661 18475 5695
rect 20806 5692 20812 5704
rect 20767 5664 20812 5692
rect 18417 5655 18475 5661
rect 20806 5652 20812 5664
rect 20864 5652 20870 5704
rect 17954 5624 17960 5636
rect 16071 5596 17960 5624
rect 16071 5593 16083 5596
rect 16025 5587 16083 5593
rect 17954 5584 17960 5596
rect 18012 5584 18018 5636
rect 18248 5624 18276 5652
rect 19613 5627 19671 5633
rect 19613 5624 19625 5627
rect 18248 5596 19625 5624
rect 19613 5593 19625 5596
rect 19659 5624 19671 5627
rect 20438 5624 20444 5636
rect 19659 5596 20444 5624
rect 19659 5593 19671 5596
rect 19613 5587 19671 5593
rect 20438 5584 20444 5596
rect 20496 5584 20502 5636
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 15672 5528 16681 5556
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 16669 5519 16727 5525
rect 18138 5516 18144 5568
rect 18196 5556 18202 5568
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 18196 5528 18245 5556
rect 18196 5516 18202 5528
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18233 5519 18291 5525
rect 18877 5559 18935 5565
rect 18877 5525 18889 5559
rect 18923 5556 18935 5559
rect 19242 5556 19248 5568
rect 18923 5528 19248 5556
rect 18923 5525 18935 5528
rect 18877 5519 18935 5525
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19705 5559 19763 5565
rect 19705 5525 19717 5559
rect 19751 5556 19763 5559
rect 19794 5556 19800 5568
rect 19751 5528 19800 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 20714 5556 20720 5568
rect 20128 5528 20720 5556
rect 20128 5516 20134 5528
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 20806 5516 20812 5568
rect 20864 5556 20870 5568
rect 20901 5559 20959 5565
rect 20901 5556 20913 5559
rect 20864 5528 20913 5556
rect 20864 5516 20870 5528
rect 20901 5525 20913 5528
rect 20947 5556 20959 5559
rect 21266 5556 21272 5568
rect 20947 5528 21272 5556
rect 20947 5525 20959 5528
rect 20901 5519 20959 5525
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 9732 5324 15853 5352
rect 9732 5312 9738 5324
rect 15841 5321 15853 5324
rect 15887 5321 15899 5355
rect 16298 5352 16304 5364
rect 16259 5324 16304 5352
rect 15841 5315 15899 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17586 5352 17592 5364
rect 17175 5324 17592 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 19797 5355 19855 5361
rect 19797 5352 19809 5355
rect 19760 5324 19809 5352
rect 19760 5312 19766 5324
rect 19797 5321 19809 5324
rect 19843 5352 19855 5355
rect 20070 5352 20076 5364
rect 19843 5324 20076 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 20165 5355 20223 5361
rect 20165 5321 20177 5355
rect 20211 5352 20223 5355
rect 20622 5352 20628 5364
rect 20211 5324 20628 5352
rect 20211 5321 20223 5324
rect 20165 5315 20223 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 15289 5287 15347 5293
rect 15289 5253 15301 5287
rect 15335 5284 15347 5287
rect 17310 5284 17316 5296
rect 15335 5256 17316 5284
rect 15335 5253 15347 5256
rect 15289 5247 15347 5253
rect 17310 5244 17316 5256
rect 17368 5244 17374 5296
rect 19242 5244 19248 5296
rect 19300 5284 19306 5296
rect 20809 5287 20867 5293
rect 20809 5284 20821 5287
rect 19300 5256 20821 5284
rect 19300 5244 19306 5256
rect 20809 5253 20821 5256
rect 20855 5253 20867 5287
rect 20809 5247 20867 5253
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17681 5219 17739 5225
rect 17681 5216 17693 5219
rect 17083 5188 17693 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17681 5185 17693 5188
rect 17727 5185 17739 5219
rect 18966 5216 18972 5228
rect 18927 5188 18972 5216
rect 17681 5179 17739 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5216 19763 5219
rect 19978 5216 19984 5228
rect 19751 5188 19984 5216
rect 19751 5185 19763 5188
rect 19705 5179 19763 5185
rect 19978 5176 19984 5188
rect 20036 5216 20042 5228
rect 20622 5216 20628 5228
rect 20036 5188 20628 5216
rect 20036 5176 20042 5188
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5117 15807 5151
rect 17310 5148 17316 5160
rect 17271 5120 17316 5148
rect 15749 5111 15807 5117
rect 15764 5080 15792 5111
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 18230 5108 18236 5160
rect 18288 5148 18294 5160
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 18288 5120 18337 5148
rect 18288 5108 18294 5120
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 18506 5108 18512 5160
rect 18564 5108 18570 5160
rect 19610 5148 19616 5160
rect 19571 5120 19616 5148
rect 19610 5108 19616 5120
rect 19668 5108 19674 5160
rect 20898 5148 20904 5160
rect 20859 5120 20904 5148
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 21082 5148 21088 5160
rect 21043 5120 21088 5148
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 18524 5080 18552 5108
rect 15764 5052 18552 5080
rect 19426 5040 19432 5092
rect 19484 5080 19490 5092
rect 19978 5080 19984 5092
rect 19484 5052 19984 5080
rect 19484 5040 19490 5052
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 20254 5040 20260 5092
rect 20312 5080 20318 5092
rect 20441 5083 20499 5089
rect 20441 5080 20453 5083
rect 20312 5052 20453 5080
rect 20312 5040 20318 5052
rect 20441 5049 20453 5052
rect 20487 5049 20499 5083
rect 20441 5043 20499 5049
rect 16390 4972 16396 5024
rect 16448 5012 16454 5024
rect 16669 5015 16727 5021
rect 16669 5012 16681 5015
rect 16448 4984 16681 5012
rect 16448 4972 16454 4984
rect 16669 4981 16681 4984
rect 16715 4981 16727 5015
rect 16669 4975 16727 4981
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 18785 5015 18843 5021
rect 18785 5012 18797 5015
rect 18564 4984 18797 5012
rect 18564 4972 18570 4984
rect 18785 4981 18797 4984
rect 18831 4981 18843 5015
rect 18785 4975 18843 4981
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 14516 4780 16957 4808
rect 14516 4768 14522 4780
rect 16945 4777 16957 4780
rect 16991 4777 17003 4811
rect 17678 4808 17684 4820
rect 16945 4771 17003 4777
rect 17052 4780 17684 4808
rect 15194 4700 15200 4752
rect 15252 4740 15258 4752
rect 16485 4743 16543 4749
rect 16485 4740 16497 4743
rect 15252 4712 16497 4740
rect 15252 4700 15258 4712
rect 16485 4709 16497 4712
rect 16531 4709 16543 4743
rect 17052 4740 17080 4780
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 19886 4808 19892 4820
rect 19484 4780 19892 4808
rect 19484 4768 19490 4780
rect 19886 4768 19892 4780
rect 19944 4808 19950 4820
rect 20162 4808 20168 4820
rect 19944 4780 20168 4808
rect 19944 4768 19950 4780
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 20346 4768 20352 4820
rect 20404 4808 20410 4820
rect 21269 4811 21327 4817
rect 21269 4808 21281 4811
rect 20404 4780 21281 4808
rect 20404 4768 20410 4780
rect 21269 4777 21281 4780
rect 21315 4777 21327 4811
rect 21269 4771 21327 4777
rect 18690 4740 18696 4752
rect 16485 4703 16543 4709
rect 16592 4712 17080 4740
rect 17144 4712 18696 4740
rect 14277 4675 14335 4681
rect 14277 4641 14289 4675
rect 14323 4672 14335 4675
rect 15930 4672 15936 4684
rect 14323 4644 15792 4672
rect 15891 4644 15936 4672
rect 14323 4641 14335 4644
rect 14277 4635 14335 4641
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6052 4576 7297 4604
rect 6052 4564 6058 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4604 14703 4607
rect 15102 4604 15108 4616
rect 14691 4576 15108 4604
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 15764 4604 15792 4644
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16592 4604 16620 4712
rect 15764 4576 16620 4604
rect 16669 4607 16727 4613
rect 15473 4567 15531 4573
rect 16669 4573 16681 4607
rect 16715 4604 16727 4607
rect 16942 4604 16948 4616
rect 16715 4576 16948 4604
rect 16715 4573 16727 4576
rect 16669 4567 16727 4573
rect 15197 4539 15255 4545
rect 15197 4505 15209 4539
rect 15243 4536 15255 4539
rect 15488 4536 15516 4567
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17144 4613 17172 4712
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 19981 4743 20039 4749
rect 19981 4709 19993 4743
rect 20027 4740 20039 4743
rect 20990 4740 20996 4752
rect 20027 4712 20996 4740
rect 20027 4709 20039 4712
rect 19981 4703 20039 4709
rect 20990 4700 20996 4712
rect 21048 4700 21054 4752
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 19518 4672 19524 4684
rect 19475 4644 19524 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4600 17647 4607
rect 17770 4604 17776 4616
rect 17696 4600 17776 4604
rect 17635 4576 17776 4600
rect 17635 4573 17724 4576
rect 17589 4572 17724 4573
rect 17589 4567 17647 4572
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 18340 4604 18368 4635
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 20530 4632 20536 4684
rect 20588 4672 20594 4684
rect 20809 4675 20867 4681
rect 20809 4672 20821 4675
rect 20588 4644 20821 4672
rect 20588 4632 20594 4644
rect 20809 4641 20821 4644
rect 20855 4641 20867 4675
rect 20809 4635 20867 4641
rect 20548 4604 20576 4632
rect 18340 4576 20576 4604
rect 17954 4536 17960 4548
rect 15243 4508 17960 4536
rect 15243 4505 15255 4508
rect 15197 4499 15255 4505
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 18509 4539 18567 4545
rect 18509 4505 18521 4539
rect 18555 4536 18567 4539
rect 19426 4536 19432 4548
rect 18555 4508 19432 4536
rect 18555 4505 18567 4508
rect 18509 4499 18567 4505
rect 19426 4496 19432 4508
rect 19484 4496 19490 4548
rect 19610 4536 19616 4548
rect 19571 4508 19616 4536
rect 19610 4496 19616 4508
rect 19668 4496 19674 4548
rect 19794 4536 19800 4548
rect 19720 4508 19800 4536
rect 7466 4468 7472 4480
rect 7427 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4468 15715 4471
rect 16298 4468 16304 4480
rect 15703 4440 16304 4468
rect 15703 4437 15715 4440
rect 15657 4431 15715 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 17405 4471 17463 4477
rect 17405 4468 17417 4471
rect 17184 4440 17417 4468
rect 17184 4428 17190 4440
rect 17405 4437 17417 4440
rect 17451 4437 17463 4471
rect 17405 4431 17463 4437
rect 17494 4428 17500 4480
rect 17552 4468 17558 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 17552 4440 18429 4468
rect 17552 4428 17558 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 18417 4431 18475 4437
rect 18877 4471 18935 4477
rect 18877 4437 18889 4471
rect 18923 4468 18935 4471
rect 19334 4468 19340 4480
rect 18923 4440 19340 4468
rect 18923 4437 18935 4440
rect 18877 4431 18935 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 19518 4468 19524 4480
rect 19479 4440 19524 4468
rect 19518 4428 19524 4440
rect 19576 4468 19582 4480
rect 19720 4468 19748 4508
rect 19794 4496 19800 4508
rect 19852 4536 19858 4548
rect 20717 4539 20775 4545
rect 20717 4536 20729 4539
rect 19852 4508 20729 4536
rect 19852 4496 19858 4508
rect 20717 4505 20729 4508
rect 20763 4505 20775 4539
rect 20717 4499 20775 4505
rect 20254 4468 20260 4480
rect 19576 4440 19748 4468
rect 20215 4440 20260 4468
rect 19576 4428 19582 4440
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 20438 4428 20444 4480
rect 20496 4468 20502 4480
rect 20625 4471 20683 4477
rect 20625 4468 20637 4471
rect 20496 4440 20637 4468
rect 20496 4428 20502 4440
rect 20625 4437 20637 4440
rect 20671 4437 20683 4471
rect 20625 4431 20683 4437
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 17034 4264 17040 4276
rect 7524 4236 17040 4264
rect 7524 4224 7530 4236
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 18230 4264 18236 4276
rect 18191 4236 18236 4264
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 19334 4264 19340 4276
rect 19295 4236 19340 4264
rect 19334 4224 19340 4236
rect 19392 4224 19398 4276
rect 19429 4267 19487 4273
rect 19429 4233 19441 4267
rect 19475 4264 19487 4267
rect 20254 4264 20260 4276
rect 19475 4236 20260 4264
rect 19475 4233 19487 4236
rect 19429 4227 19487 4233
rect 20254 4224 20260 4236
rect 20312 4224 20318 4276
rect 15102 4196 15108 4208
rect 14292 4168 15108 4196
rect 14292 4137 14320 4168
rect 15102 4156 15108 4168
rect 15160 4156 15166 4208
rect 16298 4156 16304 4208
rect 16356 4196 16362 4208
rect 19794 4196 19800 4208
rect 16356 4168 19800 4196
rect 16356 4156 16362 4168
rect 19794 4156 19800 4168
rect 19852 4196 19858 4208
rect 20806 4196 20812 4208
rect 19852 4168 20812 4196
rect 19852 4156 19858 4168
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4097 14335 4131
rect 14734 4128 14740 4140
rect 14695 4100 14740 4128
rect 14277 4091 14335 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 15378 4128 15384 4140
rect 14844 4100 15240 4128
rect 15339 4100 15384 4128
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14844 4060 14872 4100
rect 14047 4032 14872 4060
rect 15212 4060 15240 4100
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 15654 4128 15660 4140
rect 15615 4100 15660 4128
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 16114 4128 16120 4140
rect 16075 4100 16120 4128
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16816 4100 16865 4128
rect 16816 4088 16822 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17310 4128 17316 4140
rect 17175 4100 17316 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 19978 4128 19984 4140
rect 17880 4100 19656 4128
rect 19939 4100 19984 4128
rect 17880 4060 17908 4100
rect 15212 4032 17908 4060
rect 17957 4063 18015 4069
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 17957 4029 17969 4063
rect 18003 4029 18015 4063
rect 17957 4023 18015 4029
rect 16758 3952 16764 4004
rect 16816 3992 16822 4004
rect 17972 3992 18000 4023
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 18104 4032 18153 4060
rect 18104 4020 18110 4032
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 18141 4023 18199 4029
rect 18248 4032 19533 4060
rect 18248 3992 18276 4032
rect 16816 3964 17908 3992
rect 17972 3964 18276 3992
rect 18601 3995 18659 4001
rect 16816 3952 16822 3964
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14734 3924 14740 3936
rect 14507 3896 14740 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14918 3924 14924 3936
rect 14879 3896 14924 3924
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 15068 3896 15209 3924
rect 15068 3884 15074 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15197 3887 15255 3893
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16669 3927 16727 3933
rect 16669 3893 16681 3927
rect 16715 3924 16727 3927
rect 17218 3924 17224 3936
rect 16715 3896 17224 3924
rect 16715 3893 16727 3896
rect 16669 3887 16727 3893
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 17313 3927 17371 3933
rect 17313 3893 17325 3927
rect 17359 3924 17371 3927
rect 17770 3924 17776 3936
rect 17359 3896 17776 3924
rect 17359 3893 17371 3896
rect 17313 3887 17371 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 17880 3924 17908 3964
rect 18601 3961 18613 3995
rect 18647 3992 18659 3995
rect 18782 3992 18788 4004
rect 18647 3964 18788 3992
rect 18647 3961 18659 3964
rect 18601 3955 18659 3961
rect 18782 3952 18788 3964
rect 18840 3952 18846 4004
rect 18874 3952 18880 4004
rect 18932 3992 18938 4004
rect 18969 3995 19027 4001
rect 18969 3992 18981 3995
rect 18932 3964 18981 3992
rect 18932 3952 18938 3964
rect 18969 3961 18981 3964
rect 19015 3961 19027 3995
rect 18969 3955 19027 3961
rect 19058 3924 19064 3936
rect 17880 3896 19064 3924
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19352 3924 19380 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19628 4060 19656 4100
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20162 4088 20168 4140
rect 20220 4128 20226 4140
rect 20220 4100 20852 4128
rect 20220 4088 20226 4100
rect 20530 4060 20536 4072
rect 19628 4032 20536 4060
rect 19521 4023 19579 4029
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20824 4069 20852 4100
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 20162 3992 20168 4004
rect 20123 3964 20168 3992
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 22554 3924 22560 3936
rect 19352 3896 22560 3924
rect 22554 3884 22560 3896
rect 22612 3884 22618 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 16301 3723 16359 3729
rect 14792 3692 16252 3720
rect 14792 3680 14798 3692
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 14829 3655 14887 3661
rect 14829 3652 14841 3655
rect 13044 3624 14841 3652
rect 13044 3612 13050 3624
rect 14829 3621 14841 3624
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3621 15531 3655
rect 16224 3652 16252 3692
rect 16301 3689 16313 3723
rect 16347 3720 16359 3723
rect 16482 3720 16488 3732
rect 16347 3692 16488 3720
rect 16347 3689 16359 3692
rect 16301 3683 16359 3689
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 17589 3723 17647 3729
rect 17589 3720 17601 3723
rect 17368 3692 17601 3720
rect 17368 3680 17374 3692
rect 17589 3689 17601 3692
rect 17635 3689 17647 3723
rect 17589 3683 17647 3689
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 20070 3720 20076 3732
rect 18739 3692 20076 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20257 3723 20315 3729
rect 20257 3689 20269 3723
rect 20303 3720 20315 3723
rect 20898 3720 20904 3732
rect 20303 3692 20904 3720
rect 20303 3689 20315 3692
rect 20257 3683 20315 3689
rect 20898 3680 20904 3692
rect 20956 3680 20962 3732
rect 17221 3655 17279 3661
rect 16224 3624 17172 3652
rect 15473 3615 15531 3621
rect 15488 3584 15516 3615
rect 16942 3584 16948 3596
rect 13740 3556 15424 3584
rect 15488 3556 16948 3584
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13262 3448 13268 3460
rect 13223 3420 13268 3448
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 3016 3352 3065 3380
rect 3016 3340 3022 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 4338 3380 4344 3392
rect 4299 3352 4344 3380
rect 3053 3343 3111 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 13740 3389 13768 3556
rect 14366 3516 14372 3528
rect 14327 3488 14372 3516
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14734 3516 14740 3528
rect 14608 3488 14740 3516
rect 14608 3476 14614 3488
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 15010 3516 15016 3528
rect 14971 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15396 3516 15424 3556
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 17144 3584 17172 3624
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17267 3624 20944 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 20916 3596 20944 3624
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17144 3556 18061 3584
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18230 3584 18236 3596
rect 18191 3556 18236 3584
rect 18049 3547 18107 3553
rect 16022 3516 16028 3528
rect 15396 3488 16028 3516
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16390 3516 16396 3528
rect 16163 3488 16396 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3516 16819 3519
rect 16850 3516 16856 3528
rect 16807 3488 16856 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17034 3516 17040 3528
rect 16995 3488 17040 3516
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 18064 3516 18092 3547
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 19518 3584 19524 3596
rect 18524 3556 19524 3584
rect 18524 3516 18552 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 19702 3584 19708 3596
rect 19663 3556 19708 3584
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19794 3544 19800 3596
rect 19852 3584 19858 3596
rect 19852 3556 19897 3584
rect 19852 3544 19858 3556
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20772 3556 20821 3584
rect 20772 3544 20778 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 20898 3544 20904 3596
rect 20956 3544 20962 3596
rect 18064 3488 18552 3516
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 20530 3516 20536 3528
rect 18656 3488 20536 3516
rect 18656 3476 18662 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 14826 3448 14832 3460
rect 13964 3420 14832 3448
rect 13964 3408 13970 3420
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 15841 3451 15899 3457
rect 15841 3417 15853 3451
rect 15887 3448 15899 3451
rect 18782 3448 18788 3460
rect 15887 3420 18788 3448
rect 15887 3417 15899 3420
rect 15841 3411 15899 3417
rect 18782 3408 18788 3420
rect 18840 3408 18846 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 19889 3451 19947 3457
rect 19889 3448 19901 3451
rect 19576 3420 19901 3448
rect 19576 3408 19582 3420
rect 19889 3417 19901 3420
rect 19935 3417 19947 3451
rect 19889 3411 19947 3417
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3349 13783 3383
rect 14550 3380 14556 3392
rect 14511 3352 14556 3380
rect 13725 3343 13783 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 16448 3352 16589 3380
rect 16448 3340 16454 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 17954 3380 17960 3392
rect 17915 3352 17960 3380
rect 16577 3343 16635 3349
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 19978 3340 19984 3392
rect 20036 3380 20042 3392
rect 20162 3380 20168 3392
rect 20036 3352 20168 3380
rect 20036 3340 20042 3352
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 8478 3176 8484 3188
rect 2823 3148 8484 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 12529 3179 12587 3185
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12575 3148 15792 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 15562 3108 15568 3120
rect 14108 3080 15568 3108
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2556 3012 2605 3040
rect 2556 3000 2562 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3936 3012 3985 3040
rect 3936 3000 3942 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8720 3012 9045 3040
rect 8720 3000 8726 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 9033 3003 9091 3009
rect 12820 3012 13185 3040
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 12526 2904 12532 2916
rect 4203 2876 12532 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 12820 2904 12848 3012
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 13906 3040 13912 3052
rect 13679 3012 13912 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14108 3049 14136 3080
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3009 14151 3043
rect 14093 3003 14151 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14734 3040 14740 3052
rect 14599 3012 14740 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14976 3012 15209 3040
rect 14976 3000 14982 3012
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3009 15531 3043
rect 15764 3040 15792 3148
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 15896 3148 18828 3176
rect 15896 3136 15902 3148
rect 16022 3068 16028 3120
rect 16080 3108 16086 3120
rect 16080 3080 17724 3108
rect 16080 3068 16086 3080
rect 16114 3040 16120 3052
rect 15764 3012 16120 3040
rect 15473 3003 15531 3009
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 13814 2972 13820 2984
rect 12943 2944 13820 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 15488 2972 15516 3003
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3040 16267 3043
rect 16390 3040 16396 3052
rect 16255 3012 16396 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17696 3049 17724 3080
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18800 3049 18828 3148
rect 19058 3136 19064 3188
rect 19116 3176 19122 3188
rect 21174 3176 21180 3188
rect 19116 3148 21180 3176
rect 19116 3136 19122 3148
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18196 3012 18245 3040
rect 18196 3000 18202 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3009 18843 3043
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 18785 3003 18843 3009
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19886 3040 19892 3052
rect 19847 3012 19892 3040
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20680 3012 20821 3040
rect 20680 3000 20686 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 14292 2944 15516 2972
rect 14182 2904 14188 2916
rect 12820 2876 14188 2904
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 14292 2913 14320 2944
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 17402 2972 17408 2984
rect 15620 2944 17408 2972
rect 15620 2932 15626 2944
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2873 14335 2907
rect 14277 2867 14335 2873
rect 14737 2907 14795 2913
rect 14737 2873 14749 2907
rect 14783 2904 14795 2907
rect 15746 2904 15752 2916
rect 14783 2876 15752 2904
rect 14783 2873 14795 2876
rect 14737 2867 14795 2873
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 17865 2907 17923 2913
rect 17865 2873 17877 2907
rect 17911 2904 17923 2907
rect 20438 2904 20444 2916
rect 17911 2876 20444 2904
rect 17911 2873 17923 2876
rect 17865 2867 17923 2873
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 2317 2839 2375 2845
rect 2317 2805 2329 2839
rect 2363 2836 2375 2839
rect 2498 2836 2504 2848
rect 2363 2808 2504 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 3418 2836 3424 2848
rect 3375 2808 3424 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 3878 2836 3884 2848
rect 3743 2808 3884 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4798 2836 4804 2848
rect 4759 2808 4804 2836
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5258 2836 5264 2848
rect 5219 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5718 2836 5724 2848
rect 5679 2808 5724 2836
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6052 2808 6377 2836
rect 6052 2796 6058 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 6917 2839 6975 2845
rect 6917 2836 6929 2839
rect 6696 2808 6929 2836
rect 6696 2796 6702 2808
rect 6917 2805 6929 2808
rect 6963 2805 6975 2839
rect 6917 2799 6975 2805
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 7156 2808 7205 2836
rect 7156 2796 7162 2808
rect 7193 2805 7205 2808
rect 7239 2805 7251 2839
rect 7558 2836 7564 2848
rect 7519 2808 7564 2836
rect 7193 2799 7251 2805
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 8018 2836 8024 2848
rect 7979 2808 8024 2836
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 8478 2836 8484 2848
rect 8435 2808 8484 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8662 2836 8668 2848
rect 8623 2808 8668 2836
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 9456 2808 9505 2836
rect 9456 2796 9462 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9640 2808 9873 2836
rect 9640 2796 9646 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 10318 2836 10324 2848
rect 10279 2808 10324 2836
rect 9861 2799 9919 2805
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 10778 2836 10784 2848
rect 10739 2808 10784 2836
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11296 2808 11529 2836
rect 11296 2796 11302 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 13354 2836 13360 2848
rect 13315 2808 13360 2836
rect 11517 2799 11575 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 13817 2839 13875 2845
rect 13817 2805 13829 2839
rect 13863 2836 13875 2839
rect 14826 2836 14832 2848
rect 13863 2808 14832 2836
rect 13863 2805 13875 2808
rect 13817 2799 13875 2805
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 15010 2836 15016 2848
rect 14971 2808 15016 2836
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 15657 2839 15715 2845
rect 15657 2836 15669 2839
rect 15436 2808 15669 2836
rect 15436 2796 15442 2808
rect 15657 2805 15669 2808
rect 15703 2805 15715 2839
rect 16022 2836 16028 2848
rect 15983 2808 16028 2836
rect 15657 2799 15715 2805
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 16942 2836 16948 2848
rect 16903 2808 16948 2836
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18417 2839 18475 2845
rect 18417 2836 18429 2839
rect 18196 2808 18429 2836
rect 18196 2796 18202 2808
rect 18417 2805 18429 2808
rect 18463 2805 18475 2839
rect 18417 2799 18475 2805
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 18969 2839 19027 2845
rect 18969 2836 18981 2839
rect 18656 2808 18981 2836
rect 18656 2796 18662 2808
rect 18969 2805 18981 2808
rect 19015 2805 19027 2839
rect 18969 2799 19027 2805
rect 19058 2796 19064 2848
rect 19116 2836 19122 2848
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19116 2808 19533 2836
rect 19116 2796 19122 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 19521 2799 19579 2805
rect 19610 2796 19616 2848
rect 19668 2836 19674 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 19668 2808 20085 2836
rect 19668 2796 19674 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 5074 2632 5080 2644
rect 5035 2604 5080 2632
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 7282 2632 7288 2644
rect 7239 2604 7288 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 7650 2632 7656 2644
rect 7611 2604 7656 2632
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 8570 2632 8576 2644
rect 8531 2604 8576 2632
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14642 2632 14648 2644
rect 14240 2604 14648 2632
rect 14240 2592 14246 2604
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 14976 2604 15945 2632
rect 14976 2592 14982 2604
rect 15933 2601 15945 2604
rect 15979 2601 15991 2635
rect 15933 2595 15991 2601
rect 16114 2592 16120 2644
rect 16172 2632 16178 2644
rect 20530 2632 20536 2644
rect 16172 2604 20536 2632
rect 16172 2592 16178 2604
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2533 4215 2567
rect 4157 2527 4215 2533
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 8294 2564 8300 2576
rect 6043 2536 8300 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 4172 2496 4200 2527
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 9309 2567 9367 2573
rect 9309 2533 9321 2567
rect 9355 2564 9367 2567
rect 9674 2564 9680 2576
rect 9355 2536 9680 2564
rect 9355 2533 9367 2536
rect 9309 2527 9367 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 13722 2564 13728 2576
rect 11716 2536 13728 2564
rect 10686 2496 10692 2508
rect 4172 2468 10692 2496
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 2958 2428 2964 2440
rect 2823 2400 2964 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3418 2428 3424 2440
rect 3283 2400 3424 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4338 2428 4344 2440
rect 4019 2400 4344 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 4798 2428 4804 2440
rect 4479 2400 4804 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5258 2428 5264 2440
rect 4939 2400 5264 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 5718 2428 5724 2440
rect 5399 2400 5724 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 5994 2428 6000 2440
rect 5859 2400 6000 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6638 2428 6644 2440
rect 6595 2400 6644 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7098 2428 7104 2440
rect 7055 2400 7104 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7558 2428 7564 2440
rect 7515 2400 7564 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8018 2428 8024 2440
rect 7975 2400 8024 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8478 2428 8484 2440
rect 8435 2400 8484 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9398 2428 9404 2440
rect 9171 2400 9404 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9582 2428 9588 2440
rect 9543 2400 9588 2428
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10318 2428 10324 2440
rect 10091 2400 10324 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10778 2428 10784 2440
rect 10551 2400 10784 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11238 2428 11244 2440
rect 11011 2400 11244 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 2225 2363 2283 2369
rect 2225 2329 2237 2363
rect 2271 2329 2283 2363
rect 11716 2360 11744 2536
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 13998 2524 14004 2576
rect 14056 2564 14062 2576
rect 14737 2567 14795 2573
rect 14737 2564 14749 2567
rect 14056 2536 14749 2564
rect 14056 2524 14062 2536
rect 14737 2533 14749 2536
rect 14783 2533 14795 2567
rect 17126 2564 17132 2576
rect 14737 2527 14795 2533
rect 15488 2536 17132 2564
rect 15010 2496 15016 2508
rect 11900 2468 15016 2496
rect 11900 2437 11928 2468
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2397 12495 2431
rect 12986 2428 12992 2440
rect 12947 2400 12992 2428
rect 12437 2391 12495 2397
rect 2225 2323 2283 2329
rect 6748 2332 11744 2360
rect 12452 2360 12480 2391
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 14182 2428 14188 2440
rect 13587 2400 14188 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15194 2428 15200 2440
rect 14967 2400 15200 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 14274 2360 14280 2372
rect 12452 2332 14280 2360
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 2038 2292 2044 2304
rect 1903 2264 2044 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 2038 2252 2044 2264
rect 2096 2292 2102 2304
rect 2240 2292 2268 2323
rect 2096 2264 2268 2292
rect 2096 2252 2102 2264
rect 2314 2252 2320 2304
rect 2372 2292 2378 2304
rect 2961 2295 3019 2301
rect 2372 2264 2417 2292
rect 2372 2252 2378 2264
rect 2961 2261 2973 2295
rect 3007 2292 3019 2295
rect 3050 2292 3056 2304
rect 3007 2264 3056 2292
rect 3007 2261 3019 2264
rect 2961 2255 3019 2261
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 3510 2292 3516 2304
rect 3467 2264 3516 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 4614 2292 4620 2304
rect 4575 2264 4620 2292
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 5534 2292 5540 2304
rect 5495 2264 5540 2292
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 6748 2301 6776 2332
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 14384 2360 14412 2391
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15488 2437 15516 2536
rect 17126 2524 17132 2536
rect 17184 2524 17190 2576
rect 17218 2524 17224 2576
rect 17276 2564 17282 2576
rect 17957 2567 18015 2573
rect 17957 2564 17969 2567
rect 17276 2536 17969 2564
rect 17276 2524 17282 2536
rect 17957 2533 17969 2536
rect 18003 2533 18015 2567
rect 17957 2527 18015 2533
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 19981 2499 20039 2505
rect 16356 2468 17264 2496
rect 16356 2456 16362 2468
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2397 15531 2431
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15473 2391 15531 2397
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2428 16727 2431
rect 16850 2428 16856 2440
rect 16715 2400 16856 2428
rect 16715 2397 16727 2400
rect 16669 2391 16727 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17236 2437 17264 2468
rect 19981 2465 19993 2499
rect 20027 2496 20039 2499
rect 20070 2496 20076 2508
rect 20027 2468 20076 2496
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 20346 2456 20352 2508
rect 20404 2496 20410 2508
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 20404 2468 20821 2496
rect 20404 2456 20410 2468
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 20809 2459 20867 2465
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17770 2428 17776 2440
rect 17731 2400 17776 2428
rect 17221 2391 17279 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18564 2400 18613 2428
rect 18564 2388 18570 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 20254 2428 20260 2440
rect 20215 2400 20260 2428
rect 18601 2391 18659 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 20530 2428 20536 2440
rect 20443 2400 20536 2428
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 16022 2360 16028 2372
rect 14384 2332 16028 2360
rect 16022 2320 16028 2332
rect 16080 2320 16086 2372
rect 16298 2320 16304 2372
rect 16356 2360 16362 2372
rect 16356 2332 17448 2360
rect 16356 2320 16362 2332
rect 6733 2295 6791 2301
rect 6733 2261 6745 2295
rect 6779 2261 6791 2295
rect 10226 2292 10232 2304
rect 10187 2264 10232 2292
rect 6733 2255 6791 2261
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 10686 2292 10692 2304
rect 10647 2264 10692 2292
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11330 2292 11336 2304
rect 11112 2264 11336 2292
rect 11112 2252 11118 2264
rect 11330 2252 11336 2264
rect 11388 2252 11394 2304
rect 11698 2292 11704 2304
rect 11659 2264 11704 2292
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 12216 2264 12265 2292
rect 12216 2252 12222 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12253 2255 12311 2261
rect 12618 2252 12624 2304
rect 12676 2292 12682 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12676 2264 12817 2292
rect 12676 2252 12682 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13136 2264 13369 2292
rect 13136 2252 13142 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14185 2295 14243 2301
rect 14185 2292 14197 2295
rect 13596 2264 14197 2292
rect 13596 2252 13602 2264
rect 14185 2261 14197 2264
rect 14231 2261 14243 2295
rect 14185 2255 14243 2261
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14516 2264 15301 2292
rect 14516 2252 14522 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15838 2252 15844 2304
rect 15896 2292 15902 2304
rect 17420 2301 17448 2332
rect 17586 2320 17592 2372
rect 17644 2360 17650 2372
rect 20548 2360 20576 2388
rect 17644 2332 20576 2360
rect 17644 2320 17650 2332
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 15896 2264 16865 2292
rect 15896 2252 15902 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 18417 2295 18475 2301
rect 18417 2292 18429 2295
rect 17736 2264 18429 2292
rect 17736 2252 17742 2264
rect 18417 2261 18429 2264
rect 18463 2261 18475 2295
rect 18417 2255 18475 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 2314 2048 2320 2100
rect 2372 2088 2378 2100
rect 2372 2060 2774 2088
rect 2372 2048 2378 2060
rect 2746 1680 2774 2060
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 19518 2088 19524 2100
rect 10744 2060 19524 2088
rect 10744 2048 10750 2060
rect 19518 2048 19524 2060
rect 19576 2048 19582 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 11054 2020 11060 2032
rect 3108 1992 11060 2020
rect 3108 1980 3114 1992
rect 11054 1980 11060 1992
rect 11112 1980 11118 2032
rect 13814 1980 13820 2032
rect 13872 2020 13878 2032
rect 20254 2020 20260 2032
rect 13872 1992 20260 2020
rect 13872 1980 13878 1992
rect 20254 1980 20260 1992
rect 20312 1980 20318 2032
rect 4614 1912 4620 1964
rect 4672 1952 4678 1964
rect 17954 1952 17960 1964
rect 4672 1924 17960 1952
rect 4672 1912 4678 1924
rect 17954 1912 17960 1924
rect 18012 1912 18018 1964
rect 3510 1844 3516 1896
rect 3568 1884 3574 1896
rect 12342 1884 12348 1896
rect 3568 1856 12348 1884
rect 3568 1844 3574 1856
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 15102 1844 15108 1896
rect 15160 1884 15166 1896
rect 19242 1884 19248 1896
rect 15160 1856 19248 1884
rect 15160 1844 15166 1856
rect 19242 1844 19248 1856
rect 19300 1844 19306 1896
rect 5534 1776 5540 1828
rect 5592 1816 5598 1828
rect 15930 1816 15936 1828
rect 5592 1788 15936 1816
rect 5592 1776 5598 1788
rect 15930 1776 15936 1788
rect 15988 1776 15994 1828
rect 10226 1708 10232 1760
rect 10284 1748 10290 1760
rect 18046 1748 18052 1760
rect 10284 1720 18052 1748
rect 10284 1708 10290 1720
rect 18046 1708 18052 1720
rect 18104 1708 18110 1760
rect 15562 1680 15568 1692
rect 2746 1652 15568 1680
rect 15562 1640 15568 1652
rect 15620 1640 15626 1692
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 18052 20544 18104 20596
rect 7104 20476 7156 20528
rect 5724 20408 5776 20460
rect 8576 20408 8628 20460
rect 9128 20408 9180 20460
rect 11704 20408 11756 20460
rect 15292 20408 15344 20460
rect 17132 20408 17184 20460
rect 17316 20408 17368 20460
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 17592 20408 17644 20460
rect 18144 20408 18196 20460
rect 20076 20451 20128 20460
rect 8208 20340 8260 20392
rect 9496 20383 9548 20392
rect 9496 20349 9505 20383
rect 9505 20349 9539 20383
rect 9539 20349 9548 20383
rect 9496 20340 9548 20349
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 9588 20204 9640 20256
rect 10876 20204 10928 20256
rect 13176 20272 13228 20324
rect 13084 20204 13136 20256
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 20628 20408 20680 20460
rect 17960 20272 18012 20324
rect 21364 20340 21416 20392
rect 22468 20272 22520 20324
rect 15108 20247 15160 20256
rect 15108 20213 15117 20247
rect 15117 20213 15151 20247
rect 15151 20213 15160 20247
rect 15108 20204 15160 20213
rect 18052 20204 18104 20256
rect 18236 20247 18288 20256
rect 18236 20213 18245 20247
rect 18245 20213 18279 20247
rect 18279 20213 18288 20247
rect 18236 20204 18288 20213
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 18788 20204 18840 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 9128 20000 9180 20052
rect 9220 20000 9272 20052
rect 13084 20043 13136 20052
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 15108 20000 15160 20052
rect 9404 19864 9456 19916
rect 9588 19907 9640 19916
rect 9588 19873 9597 19907
rect 9597 19873 9631 19907
rect 9631 19873 9640 19907
rect 9588 19864 9640 19873
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 13176 19864 13228 19916
rect 11152 19796 11204 19848
rect 13084 19796 13136 19848
rect 17592 19932 17644 19984
rect 11244 19728 11296 19780
rect 15292 19796 15344 19848
rect 17500 19864 17552 19916
rect 21364 19907 21416 19916
rect 16856 19796 16908 19848
rect 7748 19660 7800 19712
rect 8668 19660 8720 19712
rect 10508 19660 10560 19712
rect 12624 19660 12676 19712
rect 14924 19703 14976 19712
rect 14924 19669 14933 19703
rect 14933 19669 14967 19703
rect 14967 19669 14976 19703
rect 14924 19660 14976 19669
rect 16396 19660 16448 19712
rect 21364 19873 21373 19907
rect 21373 19873 21407 19907
rect 21407 19873 21416 19907
rect 21364 19864 21416 19873
rect 19708 19728 19760 19780
rect 21548 19728 21600 19780
rect 17592 19660 17644 19712
rect 19616 19703 19668 19712
rect 19616 19669 19625 19703
rect 19625 19669 19659 19703
rect 19659 19669 19668 19703
rect 19616 19660 19668 19669
rect 20812 19660 20864 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 7104 19499 7156 19508
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 9496 19456 9548 19508
rect 10508 19456 10560 19508
rect 11980 19456 12032 19508
rect 8852 19431 8904 19440
rect 8852 19397 8861 19431
rect 8861 19397 8895 19431
rect 8895 19397 8904 19431
rect 8852 19388 8904 19397
rect 9864 19388 9916 19440
rect 10784 19388 10836 19440
rect 10876 19431 10928 19440
rect 10876 19397 10894 19431
rect 10894 19397 10928 19431
rect 10876 19388 10928 19397
rect 11060 19388 11112 19440
rect 14924 19456 14976 19508
rect 18144 19456 18196 19508
rect 18512 19456 18564 19508
rect 18880 19456 18932 19508
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 9404 19320 9456 19372
rect 16396 19388 16448 19440
rect 8024 19295 8076 19304
rect 8024 19261 8033 19295
rect 8033 19261 8067 19295
rect 8067 19261 8076 19295
rect 8024 19252 8076 19261
rect 11152 19295 11204 19304
rect 9864 19184 9916 19236
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 11152 19261 11161 19295
rect 11161 19261 11195 19295
rect 11195 19261 11204 19295
rect 11152 19252 11204 19261
rect 10508 19116 10560 19168
rect 11244 19116 11296 19168
rect 13820 19116 13872 19168
rect 15936 19252 15988 19304
rect 18052 19320 18104 19372
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 17960 19116 18012 19168
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 20628 19116 20680 19168
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 8024 18912 8076 18964
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 11704 18912 11756 18964
rect 16304 18912 16356 18964
rect 11888 18844 11940 18896
rect 8392 18708 8444 18760
rect 11152 18708 11204 18760
rect 9496 18640 9548 18692
rect 8392 18615 8444 18624
rect 8392 18581 8401 18615
rect 8401 18581 8435 18615
rect 8435 18581 8444 18615
rect 8392 18572 8444 18581
rect 9220 18572 9272 18624
rect 12624 18683 12676 18692
rect 12624 18649 12642 18683
rect 12642 18649 12676 18683
rect 12624 18640 12676 18649
rect 13820 18708 13872 18760
rect 17592 18776 17644 18828
rect 18696 18751 18748 18760
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 17132 18640 17184 18692
rect 15936 18615 15988 18624
rect 15936 18581 15945 18615
rect 15945 18581 15979 18615
rect 15979 18581 15988 18615
rect 15936 18572 15988 18581
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 22376 18708 22428 18760
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 20352 18640 20404 18692
rect 17960 18572 18012 18581
rect 19156 18572 19208 18624
rect 19892 18572 19944 18624
rect 20720 18572 20772 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 8576 18368 8628 18420
rect 9220 18411 9272 18420
rect 9220 18377 9229 18411
rect 9229 18377 9263 18411
rect 9263 18377 9272 18411
rect 9220 18368 9272 18377
rect 11152 18368 11204 18420
rect 11704 18368 11756 18420
rect 11888 18368 11940 18420
rect 17316 18368 17368 18420
rect 8392 18300 8444 18352
rect 16948 18300 17000 18352
rect 13176 18275 13228 18284
rect 13176 18241 13194 18275
rect 13194 18241 13228 18275
rect 13176 18232 13228 18241
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 9496 18164 9548 18173
rect 13268 18028 13320 18080
rect 16764 18232 16816 18284
rect 17500 18232 17552 18284
rect 19156 18275 19208 18284
rect 19156 18241 19165 18275
rect 19165 18241 19199 18275
rect 19199 18241 19208 18275
rect 19156 18232 19208 18241
rect 19524 18232 19576 18284
rect 20260 18275 20312 18284
rect 20260 18241 20294 18275
rect 20294 18241 20312 18275
rect 20260 18232 20312 18241
rect 16304 18207 16356 18216
rect 16304 18173 16313 18207
rect 16313 18173 16347 18207
rect 16347 18173 16356 18207
rect 16304 18164 16356 18173
rect 17960 18096 18012 18148
rect 19616 18139 19668 18148
rect 19616 18105 19625 18139
rect 19625 18105 19659 18139
rect 19659 18105 19668 18139
rect 19616 18096 19668 18105
rect 18052 18028 18104 18080
rect 21548 18028 21600 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 18880 17867 18932 17876
rect 18880 17833 18889 17867
rect 18889 17833 18923 17867
rect 18923 17833 18932 17867
rect 18880 17824 18932 17833
rect 15568 17756 15620 17808
rect 20720 17824 20772 17876
rect 11888 17620 11940 17672
rect 17960 17620 18012 17672
rect 18604 17620 18656 17672
rect 19248 17620 19300 17672
rect 21180 17620 21232 17672
rect 19892 17552 19944 17604
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 13268 17484 13320 17536
rect 15844 17484 15896 17536
rect 16304 17484 16356 17536
rect 19708 17484 19760 17536
rect 20260 17484 20312 17536
rect 20536 17484 20588 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 15844 17212 15896 17264
rect 17960 17212 18012 17264
rect 13728 17144 13780 17196
rect 15568 17144 15620 17196
rect 18512 17144 18564 17196
rect 20444 17212 20496 17264
rect 19708 17187 19760 17196
rect 19708 17153 19742 17187
rect 19742 17153 19760 17187
rect 21088 17187 21140 17196
rect 13268 17008 13320 17060
rect 19708 17144 19760 17153
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 19248 17076 19300 17128
rect 17316 17008 17368 17060
rect 18972 17051 19024 17060
rect 18972 17017 18981 17051
rect 18981 17017 19015 17051
rect 19015 17017 19024 17051
rect 18972 17008 19024 17017
rect 20628 17008 20680 17060
rect 14556 16940 14608 16992
rect 17684 16940 17736 16992
rect 20720 16940 20772 16992
rect 22744 16940 22796 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 10508 16779 10560 16788
rect 10508 16745 10517 16779
rect 10517 16745 10551 16779
rect 10551 16745 10560 16779
rect 10508 16736 10560 16745
rect 11704 16736 11756 16788
rect 9404 16643 9456 16652
rect 9404 16609 9413 16643
rect 9413 16609 9447 16643
rect 9447 16609 9456 16643
rect 9404 16600 9456 16609
rect 9864 16600 9916 16652
rect 18512 16736 18564 16788
rect 18788 16736 18840 16788
rect 13268 16600 13320 16652
rect 11796 16532 11848 16584
rect 15844 16532 15896 16584
rect 17960 16575 18012 16584
rect 17960 16541 17969 16575
rect 17969 16541 18003 16575
rect 18003 16541 18012 16575
rect 17960 16532 18012 16541
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 8668 16396 8720 16448
rect 10968 16396 11020 16448
rect 14556 16507 14608 16516
rect 14556 16473 14590 16507
rect 14590 16473 14608 16507
rect 14556 16464 14608 16473
rect 16212 16507 16264 16516
rect 13728 16396 13780 16448
rect 16212 16473 16246 16507
rect 16246 16473 16264 16507
rect 16212 16464 16264 16473
rect 17868 16464 17920 16516
rect 19248 16532 19300 16584
rect 22192 16532 22244 16584
rect 17500 16396 17552 16448
rect 19524 16464 19576 16516
rect 20812 16464 20864 16516
rect 22100 16464 22152 16516
rect 20076 16396 20128 16448
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 19156 16192 19208 16244
rect 9588 16056 9640 16108
rect 17960 16056 18012 16108
rect 20720 16124 20772 16176
rect 19800 16056 19852 16108
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 19248 15988 19300 16040
rect 9864 15852 9916 15904
rect 10968 15852 11020 15904
rect 13268 15895 13320 15904
rect 13268 15861 13277 15895
rect 13277 15861 13311 15895
rect 13311 15861 13320 15895
rect 13268 15852 13320 15861
rect 16948 15852 17000 15904
rect 17408 15852 17460 15904
rect 20996 15852 21048 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 15844 15555 15896 15564
rect 15844 15521 15853 15555
rect 15853 15521 15887 15555
rect 15887 15521 15896 15555
rect 15844 15512 15896 15521
rect 16304 15512 16356 15564
rect 18052 15512 18104 15564
rect 21640 15648 21692 15700
rect 12072 15376 12124 15428
rect 9588 15308 9640 15360
rect 20628 15444 20680 15496
rect 18236 15376 18288 15428
rect 13268 15308 13320 15360
rect 14832 15308 14884 15360
rect 19248 15308 19300 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 21364 15308 21416 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 18328 15104 18380 15156
rect 13820 14968 13872 15020
rect 14832 15011 14884 15020
rect 14832 14977 14866 15011
rect 14866 14977 14884 15011
rect 14832 14968 14884 14977
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 20628 15036 20680 15088
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 20812 14968 20864 15020
rect 21456 14900 21508 14952
rect 12072 14764 12124 14816
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 18144 14764 18196 14816
rect 18236 14764 18288 14816
rect 18972 14764 19024 14816
rect 19800 14764 19852 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 14832 14560 14884 14612
rect 18052 14560 18104 14612
rect 19524 14603 19576 14612
rect 19524 14569 19533 14603
rect 19533 14569 19567 14603
rect 19567 14569 19576 14603
rect 19524 14560 19576 14569
rect 11980 14356 12032 14408
rect 13636 14356 13688 14408
rect 11704 14220 11756 14272
rect 15936 14356 15988 14408
rect 16304 14356 16356 14408
rect 18512 14356 18564 14408
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 20628 14356 20680 14408
rect 16948 14288 17000 14340
rect 17224 14331 17276 14340
rect 17224 14297 17253 14331
rect 17253 14297 17276 14331
rect 17224 14288 17276 14297
rect 20996 14288 21048 14340
rect 12900 14220 12952 14272
rect 18328 14220 18380 14272
rect 20812 14220 20864 14272
rect 22652 14220 22704 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 10048 14016 10100 14068
rect 13820 14016 13872 14068
rect 16948 14016 17000 14068
rect 17684 14016 17736 14068
rect 18420 14016 18472 14068
rect 19616 14016 19668 14068
rect 20720 14059 20772 14068
rect 9404 13948 9456 14000
rect 15752 13948 15804 14000
rect 17224 13948 17276 14000
rect 18880 13948 18932 14000
rect 19984 13948 20036 14000
rect 20720 14025 20729 14059
rect 20729 14025 20763 14059
rect 20763 14025 20772 14059
rect 20720 14016 20772 14025
rect 21456 13948 21508 14000
rect 22284 13948 22336 14000
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 12808 13880 12860 13932
rect 16304 13880 16356 13932
rect 18512 13923 18564 13932
rect 18512 13889 18521 13923
rect 18521 13889 18555 13923
rect 18555 13889 18564 13923
rect 18512 13880 18564 13889
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 20996 13880 21048 13932
rect 11980 13855 12032 13864
rect 9588 13744 9640 13796
rect 11152 13676 11204 13728
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 20628 13812 20680 13864
rect 21456 13812 21508 13864
rect 13636 13719 13688 13728
rect 13636 13685 13645 13719
rect 13645 13685 13679 13719
rect 13679 13685 13688 13719
rect 13636 13676 13688 13685
rect 17132 13676 17184 13728
rect 17500 13676 17552 13728
rect 19984 13676 20036 13728
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 21364 13515 21416 13524
rect 21364 13481 21373 13515
rect 21373 13481 21407 13515
rect 21407 13481 21416 13515
rect 21364 13472 21416 13481
rect 22560 13472 22612 13524
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 14556 13336 14608 13388
rect 18512 13336 18564 13388
rect 19984 13379 20036 13388
rect 19984 13345 19993 13379
rect 19993 13345 20027 13379
rect 20027 13345 20036 13379
rect 19984 13336 20036 13345
rect 13636 13268 13688 13320
rect 16028 13268 16080 13320
rect 16120 13268 16172 13320
rect 20076 13268 20128 13320
rect 11704 13200 11756 13252
rect 12808 13132 12860 13184
rect 16212 13132 16264 13184
rect 17960 13200 18012 13252
rect 18144 13243 18196 13252
rect 18144 13209 18162 13243
rect 18162 13209 18196 13243
rect 18144 13200 18196 13209
rect 20352 13200 20404 13252
rect 16396 13132 16448 13184
rect 17224 13132 17276 13184
rect 20720 13132 20772 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 16120 12928 16172 12980
rect 18696 12971 18748 12980
rect 18696 12937 18705 12971
rect 18705 12937 18739 12971
rect 18739 12937 18748 12971
rect 18696 12928 18748 12937
rect 21088 12928 21140 12980
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 18972 12860 19024 12912
rect 20628 12835 20680 12844
rect 12072 12724 12124 12776
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 15292 12724 15344 12776
rect 17592 12767 17644 12776
rect 14740 12656 14792 12708
rect 13176 12588 13228 12640
rect 16948 12588 17000 12640
rect 17592 12733 17601 12767
rect 17601 12733 17635 12767
rect 17635 12733 17644 12767
rect 17592 12724 17644 12733
rect 19892 12724 19944 12776
rect 19064 12656 19116 12708
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 20904 12792 20956 12844
rect 20812 12656 20864 12708
rect 21088 12656 21140 12708
rect 21364 12588 21416 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 11888 12384 11940 12436
rect 15016 12384 15068 12436
rect 13636 12316 13688 12368
rect 13728 12316 13780 12368
rect 16212 12384 16264 12436
rect 18972 12384 19024 12436
rect 19708 12384 19760 12436
rect 21272 12427 21324 12436
rect 21272 12393 21281 12427
rect 21281 12393 21315 12427
rect 21315 12393 21324 12427
rect 21272 12384 21324 12393
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 11244 12248 11296 12300
rect 13268 12248 13320 12300
rect 13820 12248 13872 12300
rect 15844 12291 15896 12300
rect 15844 12257 15853 12291
rect 15853 12257 15887 12291
rect 15887 12257 15896 12291
rect 15844 12248 15896 12257
rect 16948 12316 17000 12368
rect 17500 12316 17552 12368
rect 17040 12248 17092 12300
rect 7840 12180 7892 12232
rect 15476 12180 15528 12232
rect 16396 12180 16448 12232
rect 11244 12044 11296 12096
rect 13820 12112 13872 12164
rect 17960 12180 18012 12232
rect 20904 12316 20956 12368
rect 21088 12316 21140 12368
rect 20260 12248 20312 12300
rect 13176 12044 13228 12096
rect 15200 12044 15252 12096
rect 15384 12044 15436 12096
rect 16028 12044 16080 12096
rect 19524 12112 19576 12164
rect 20076 12180 20128 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 17500 12044 17552 12096
rect 18420 12044 18472 12096
rect 18604 12044 18656 12096
rect 19800 12044 19852 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 9312 11840 9364 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 15476 11840 15528 11892
rect 17592 11840 17644 11892
rect 19064 11840 19116 11892
rect 19524 11840 19576 11892
rect 19708 11883 19760 11892
rect 19708 11849 19717 11883
rect 19717 11849 19751 11883
rect 19751 11849 19760 11883
rect 19708 11840 19760 11849
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12624 11679 12676 11688
rect 12440 11636 12492 11645
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 13636 11772 13688 11824
rect 15660 11704 15712 11756
rect 18052 11704 18104 11756
rect 19616 11747 19668 11756
rect 12808 11636 12860 11688
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 17684 11636 17736 11688
rect 16948 11568 17000 11620
rect 17500 11568 17552 11620
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 21456 11840 21508 11892
rect 20720 11772 20772 11824
rect 18788 11679 18840 11688
rect 18788 11645 18797 11679
rect 18797 11645 18831 11679
rect 18831 11645 18840 11679
rect 18788 11636 18840 11645
rect 19984 11636 20036 11688
rect 21272 11636 21324 11688
rect 20444 11568 20496 11620
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 16028 11500 16080 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 17040 11500 17092 11552
rect 19524 11500 19576 11552
rect 22192 11500 22244 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 14832 11296 14884 11348
rect 17684 11296 17736 11348
rect 17868 11296 17920 11348
rect 18420 11296 18472 11348
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 19984 11296 20036 11348
rect 21180 11339 21232 11348
rect 12440 11228 12492 11280
rect 11704 11160 11756 11212
rect 16856 11228 16908 11280
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 15844 11160 15896 11212
rect 18052 11203 18104 11212
rect 17592 11135 17644 11144
rect 7288 11024 7340 11076
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 19064 11160 19116 11212
rect 19340 11135 19392 11144
rect 17960 11024 18012 11076
rect 19340 11101 19349 11135
rect 19349 11101 19383 11135
rect 19383 11101 19392 11135
rect 19340 11092 19392 11101
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20260 11092 20312 11144
rect 21640 11228 21692 11280
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 21456 11024 21508 11076
rect 15292 10999 15344 11008
rect 15292 10965 15301 10999
rect 15301 10965 15335 10999
rect 15335 10965 15344 10999
rect 15292 10956 15344 10965
rect 16948 10956 17000 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 15292 10752 15344 10804
rect 15660 10752 15712 10804
rect 17316 10752 17368 10804
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 18512 10752 18564 10804
rect 19340 10752 19392 10804
rect 20536 10795 20588 10804
rect 17868 10684 17920 10736
rect 20536 10761 20545 10795
rect 20545 10761 20579 10795
rect 20579 10761 20588 10795
rect 20536 10752 20588 10761
rect 20812 10752 20864 10804
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 21456 10752 21508 10804
rect 18696 10616 18748 10668
rect 19892 10659 19944 10668
rect 15016 10548 15068 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 18604 10548 18656 10600
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 17960 10480 18012 10532
rect 20628 10480 20680 10532
rect 15936 10412 15988 10464
rect 19524 10412 19576 10464
rect 22376 10412 22428 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 17592 10208 17644 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 20812 10208 20864 10260
rect 11152 10140 11204 10192
rect 15936 10140 15988 10192
rect 17224 10140 17276 10192
rect 20076 10183 20128 10192
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 17408 10072 17460 10124
rect 20076 10149 20085 10183
rect 20085 10149 20119 10183
rect 20119 10149 20128 10183
rect 20076 10140 20128 10149
rect 15200 10004 15252 10056
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 16948 10004 17000 10056
rect 17500 10004 17552 10056
rect 18236 10004 18288 10056
rect 22744 10072 22796 10124
rect 8116 9936 8168 9988
rect 17224 9936 17276 9988
rect 20168 9936 20220 9988
rect 15200 9868 15252 9920
rect 16948 9868 17000 9920
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 20720 9911 20772 9920
rect 18328 9868 18380 9877
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 20996 9868 21048 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 17500 9707 17552 9716
rect 17500 9673 17509 9707
rect 17509 9673 17543 9707
rect 17543 9673 17552 9707
rect 17500 9664 17552 9673
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 11796 9596 11848 9648
rect 15200 9639 15252 9648
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 15200 9605 15209 9639
rect 15209 9605 15243 9639
rect 15243 9605 15252 9639
rect 15200 9596 15252 9605
rect 19892 9664 19944 9716
rect 20168 9707 20220 9716
rect 20168 9673 20177 9707
rect 20177 9673 20211 9707
rect 20211 9673 20220 9707
rect 20168 9664 20220 9673
rect 19616 9596 19668 9648
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 18236 9528 18288 9580
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 12164 9435 12216 9444
rect 12164 9401 12173 9435
rect 12173 9401 12207 9435
rect 12207 9401 12216 9435
rect 12164 9392 12216 9401
rect 12900 9460 12952 9512
rect 15568 9460 15620 9512
rect 18420 9460 18472 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 20904 9460 20956 9512
rect 15016 9392 15068 9444
rect 17868 9392 17920 9444
rect 20352 9392 20404 9444
rect 21640 9528 21692 9580
rect 21180 9367 21232 9376
rect 21180 9333 21189 9367
rect 21189 9333 21223 9367
rect 21223 9333 21232 9367
rect 21180 9324 21232 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 15568 9163 15620 9172
rect 15568 9129 15577 9163
rect 15577 9129 15611 9163
rect 15611 9129 15620 9163
rect 15568 9120 15620 9129
rect 17316 9120 17368 9172
rect 18328 9120 18380 9172
rect 19984 9120 20036 9172
rect 20628 9120 20680 9172
rect 21088 9163 21140 9172
rect 21088 9129 21097 9163
rect 21097 9129 21131 9163
rect 21131 9129 21140 9163
rect 21088 9120 21140 9129
rect 15844 9052 15896 9104
rect 16120 8984 16172 9036
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 18420 8984 18472 9036
rect 5080 8780 5132 8832
rect 7656 8780 7708 8832
rect 18328 8916 18380 8968
rect 18972 8916 19024 8968
rect 15016 8780 15068 8832
rect 19708 8916 19760 8968
rect 19892 8984 19944 9036
rect 20904 8984 20956 9036
rect 20628 8848 20680 8900
rect 17132 8780 17184 8832
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 18052 8780 18104 8832
rect 19340 8780 19392 8832
rect 19616 8780 19668 8832
rect 20352 8823 20404 8832
rect 20352 8789 20361 8823
rect 20361 8789 20395 8823
rect 20395 8789 20404 8823
rect 20352 8780 20404 8789
rect 20812 8780 20864 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 17960 8619 18012 8628
rect 9220 8508 9272 8560
rect 17500 8508 17552 8560
rect 17960 8585 17969 8619
rect 17969 8585 18003 8619
rect 18003 8585 18012 8619
rect 17960 8576 18012 8585
rect 19340 8576 19392 8628
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 20720 8619 20772 8628
rect 20720 8585 20729 8619
rect 20729 8585 20763 8619
rect 20763 8585 20772 8619
rect 20720 8576 20772 8585
rect 21272 8576 21324 8628
rect 17132 8440 17184 8492
rect 17960 8440 18012 8492
rect 18236 8440 18288 8492
rect 16304 8372 16356 8424
rect 16120 8304 16172 8356
rect 18788 8440 18840 8492
rect 19248 8440 19300 8492
rect 20260 8508 20312 8560
rect 21364 8483 21416 8492
rect 21364 8449 21373 8483
rect 21373 8449 21407 8483
rect 21407 8449 21416 8483
rect 21364 8440 21416 8449
rect 20168 8415 20220 8424
rect 18696 8304 18748 8356
rect 20168 8381 20177 8415
rect 20177 8381 20211 8415
rect 20211 8381 20220 8415
rect 20168 8372 20220 8381
rect 22100 8372 22152 8424
rect 21272 8304 21324 8356
rect 15476 8236 15528 8288
rect 19892 8236 19944 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 17776 8032 17828 8084
rect 18788 8032 18840 8084
rect 20352 8075 20404 8084
rect 20352 8041 20361 8075
rect 20361 8041 20395 8075
rect 20395 8041 20404 8075
rect 20352 8032 20404 8041
rect 18696 7964 18748 8016
rect 21180 7964 21232 8016
rect 18144 7896 18196 7948
rect 19616 7896 19668 7948
rect 20076 7896 20128 7948
rect 20720 7896 20772 7948
rect 22284 7896 22336 7948
rect 18972 7828 19024 7880
rect 16304 7760 16356 7812
rect 19708 7828 19760 7880
rect 22468 7828 22520 7880
rect 18144 7735 18196 7744
rect 18144 7701 18153 7735
rect 18153 7701 18187 7735
rect 18187 7701 18196 7735
rect 18144 7692 18196 7701
rect 18420 7692 18472 7744
rect 19892 7692 19944 7744
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 15752 7488 15804 7540
rect 17868 7488 17920 7540
rect 19524 7488 19576 7540
rect 19708 7488 19760 7540
rect 20812 7488 20864 7540
rect 15292 7420 15344 7472
rect 18420 7420 18472 7472
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 15568 7284 15620 7336
rect 18052 7284 18104 7336
rect 18880 7420 18932 7472
rect 19064 7420 19116 7472
rect 18788 7352 18840 7404
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 20628 7352 20680 7404
rect 21456 7352 21508 7404
rect 20720 7216 20772 7268
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 18052 7148 18104 7200
rect 21180 7191 21232 7200
rect 21180 7157 21189 7191
rect 21189 7157 21223 7191
rect 21223 7157 21232 7191
rect 21180 7148 21232 7157
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 19432 6944 19484 6996
rect 19892 6944 19944 6996
rect 17316 6808 17368 6860
rect 17592 6808 17644 6860
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 18604 6876 18656 6928
rect 19984 6876 20036 6928
rect 20628 6876 20680 6928
rect 19524 6808 19576 6860
rect 19800 6808 19852 6860
rect 17500 6740 17552 6792
rect 18328 6740 18380 6792
rect 18972 6740 19024 6792
rect 17408 6604 17460 6656
rect 17592 6647 17644 6656
rect 17592 6613 17601 6647
rect 17601 6613 17635 6647
rect 17635 6613 17644 6647
rect 17592 6604 17644 6613
rect 17776 6604 17828 6656
rect 19524 6672 19576 6724
rect 18972 6604 19024 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 20076 6808 20128 6860
rect 21088 6808 21140 6860
rect 21548 6808 21600 6860
rect 19892 6672 19944 6724
rect 21364 6715 21416 6724
rect 20076 6604 20128 6656
rect 20168 6604 20220 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 21364 6681 21373 6715
rect 21373 6681 21407 6715
rect 21407 6681 21416 6715
rect 21364 6672 21416 6681
rect 22652 6604 22704 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 18144 6443 18196 6452
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 19248 6400 19300 6452
rect 20536 6400 20588 6452
rect 18052 6332 18104 6384
rect 17500 6264 17552 6316
rect 17776 6264 17828 6316
rect 17960 6264 18012 6316
rect 18512 6264 18564 6316
rect 18604 6239 18656 6248
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 20352 6264 20404 6316
rect 20444 6196 20496 6248
rect 20904 6239 20956 6248
rect 20904 6205 20913 6239
rect 20913 6205 20947 6239
rect 20947 6205 20956 6239
rect 20904 6196 20956 6205
rect 10692 6128 10744 6180
rect 13176 6128 13228 6180
rect 15660 6128 15712 6180
rect 14832 6060 14884 6112
rect 17776 6060 17828 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 14648 5856 14700 5908
rect 18604 5856 18656 5908
rect 20444 5899 20496 5908
rect 20444 5865 20453 5899
rect 20453 5865 20487 5899
rect 20487 5865 20496 5899
rect 20444 5856 20496 5865
rect 14372 5788 14424 5840
rect 15752 5720 15804 5772
rect 17868 5788 17920 5840
rect 17408 5720 17460 5772
rect 19892 5763 19944 5772
rect 14280 5584 14332 5636
rect 17684 5652 17736 5704
rect 18236 5652 18288 5704
rect 19892 5729 19901 5763
rect 19901 5729 19935 5763
rect 19935 5729 19944 5763
rect 19892 5720 19944 5729
rect 20720 5720 20772 5772
rect 20812 5695 20864 5704
rect 20812 5661 20821 5695
rect 20821 5661 20855 5695
rect 20855 5661 20864 5695
rect 20812 5652 20864 5661
rect 17960 5584 18012 5636
rect 20444 5584 20496 5636
rect 18144 5516 18196 5568
rect 19248 5516 19300 5568
rect 19800 5516 19852 5568
rect 20076 5516 20128 5568
rect 20720 5516 20772 5568
rect 20812 5516 20864 5568
rect 21272 5516 21324 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 9680 5312 9732 5364
rect 16304 5355 16356 5364
rect 16304 5321 16313 5355
rect 16313 5321 16347 5355
rect 16347 5321 16356 5355
rect 16304 5312 16356 5321
rect 17592 5312 17644 5364
rect 19708 5312 19760 5364
rect 20076 5312 20128 5364
rect 20628 5312 20680 5364
rect 17316 5244 17368 5296
rect 19248 5244 19300 5296
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 19984 5176 20036 5228
rect 20628 5176 20680 5228
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 18236 5108 18288 5160
rect 18512 5108 18564 5160
rect 19616 5151 19668 5160
rect 19616 5117 19625 5151
rect 19625 5117 19659 5151
rect 19659 5117 19668 5151
rect 19616 5108 19668 5117
rect 20904 5151 20956 5160
rect 20904 5117 20913 5151
rect 20913 5117 20947 5151
rect 20947 5117 20956 5151
rect 20904 5108 20956 5117
rect 21088 5151 21140 5160
rect 21088 5117 21097 5151
rect 21097 5117 21131 5151
rect 21131 5117 21140 5151
rect 21088 5108 21140 5117
rect 19432 5040 19484 5092
rect 19984 5040 20036 5092
rect 20260 5040 20312 5092
rect 16396 4972 16448 5024
rect 18512 4972 18564 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 14464 4768 14516 4820
rect 15200 4700 15252 4752
rect 17684 4768 17736 4820
rect 19432 4768 19484 4820
rect 19892 4768 19944 4820
rect 20168 4768 20220 4820
rect 20352 4768 20404 4820
rect 15936 4675 15988 4684
rect 6000 4564 6052 4616
rect 15108 4564 15160 4616
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16948 4564 17000 4616
rect 18696 4700 18748 4752
rect 20996 4700 21048 4752
rect 17776 4564 17828 4616
rect 19524 4632 19576 4684
rect 20536 4632 20588 4684
rect 17960 4496 18012 4548
rect 19432 4496 19484 4548
rect 19616 4539 19668 4548
rect 19616 4505 19625 4539
rect 19625 4505 19659 4539
rect 19659 4505 19668 4539
rect 19616 4496 19668 4505
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 16304 4428 16356 4480
rect 17132 4428 17184 4480
rect 17500 4428 17552 4480
rect 19340 4428 19392 4480
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19800 4496 19852 4548
rect 20260 4471 20312 4480
rect 19524 4428 19576 4437
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20444 4428 20496 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 7472 4224 7524 4276
rect 17040 4224 17092 4276
rect 18236 4267 18288 4276
rect 18236 4233 18245 4267
rect 18245 4233 18279 4267
rect 18279 4233 18288 4267
rect 18236 4224 18288 4233
rect 19340 4267 19392 4276
rect 19340 4233 19349 4267
rect 19349 4233 19383 4267
rect 19383 4233 19392 4267
rect 19340 4224 19392 4233
rect 20260 4224 20312 4276
rect 15108 4156 15160 4208
rect 16304 4156 16356 4208
rect 19800 4156 19852 4208
rect 20812 4156 20864 4208
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16764 4088 16816 4140
rect 17316 4088 17368 4140
rect 19984 4131 20036 4140
rect 16764 3952 16816 4004
rect 18052 4020 18104 4072
rect 14740 3884 14792 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 15016 3884 15068 3936
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 17224 3884 17276 3936
rect 17776 3884 17828 3936
rect 18788 3952 18840 4004
rect 18880 3952 18932 4004
rect 19064 3884 19116 3936
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 20168 4088 20220 4140
rect 20536 4063 20588 4072
rect 20536 4029 20545 4063
rect 20545 4029 20579 4063
rect 20579 4029 20588 4063
rect 20536 4020 20588 4029
rect 20168 3995 20220 4004
rect 20168 3961 20177 3995
rect 20177 3961 20211 3995
rect 20211 3961 20220 3995
rect 20168 3952 20220 3961
rect 22560 3884 22612 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 14740 3680 14792 3732
rect 12992 3612 13044 3664
rect 16488 3680 16540 3732
rect 17316 3680 17368 3732
rect 20076 3680 20128 3732
rect 20904 3680 20956 3732
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 13268 3451 13320 3460
rect 13268 3417 13277 3451
rect 13277 3417 13311 3451
rect 13311 3417 13320 3451
rect 13268 3408 13320 3417
rect 2964 3340 3016 3392
rect 4344 3383 4396 3392
rect 4344 3349 4353 3383
rect 4353 3349 4387 3383
rect 4387 3349 4396 3383
rect 4344 3340 4396 3349
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 14556 3476 14608 3528
rect 14740 3476 14792 3528
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 16948 3544 17000 3596
rect 18236 3587 18288 3596
rect 16028 3476 16080 3528
rect 16396 3476 16448 3528
rect 16856 3476 16908 3528
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 18236 3553 18245 3587
rect 18245 3553 18279 3587
rect 18279 3553 18288 3587
rect 18236 3544 18288 3553
rect 19524 3544 19576 3596
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 20720 3544 20772 3596
rect 20904 3544 20956 3596
rect 18604 3476 18656 3528
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 13912 3408 13964 3460
rect 14832 3408 14884 3460
rect 18788 3451 18840 3460
rect 18788 3417 18797 3451
rect 18797 3417 18831 3451
rect 18831 3417 18840 3451
rect 18788 3408 18840 3417
rect 19524 3408 19576 3460
rect 14556 3383 14608 3392
rect 14556 3349 14565 3383
rect 14565 3349 14599 3383
rect 14599 3349 14608 3383
rect 14556 3340 14608 3349
rect 16396 3340 16448 3392
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 19984 3340 20036 3392
rect 20168 3340 20220 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 8484 3136 8536 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 2504 3000 2556 3052
rect 3884 3000 3936 3052
rect 8668 3000 8720 3052
rect 12532 2864 12584 2916
rect 13912 3000 13964 3052
rect 15568 3068 15620 3120
rect 14740 3000 14792 3052
rect 14924 3000 14976 3052
rect 15844 3136 15896 3188
rect 16028 3068 16080 3120
rect 13820 2932 13872 2984
rect 16120 3000 16172 3052
rect 16396 3000 16448 3052
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 18144 3000 18196 3052
rect 19064 3136 19116 3188
rect 21180 3136 21232 3188
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 19892 3043 19944 3052
rect 19892 3009 19901 3043
rect 19901 3009 19935 3043
rect 19935 3009 19944 3043
rect 19892 3000 19944 3009
rect 20628 3000 20680 3052
rect 14188 2864 14240 2916
rect 15568 2932 15620 2984
rect 17408 2932 17460 2984
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 15752 2864 15804 2916
rect 20444 2864 20496 2916
rect 2504 2796 2556 2848
rect 3424 2796 3476 2848
rect 3884 2796 3936 2848
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 5724 2839 5776 2848
rect 5724 2805 5733 2839
rect 5733 2805 5767 2839
rect 5767 2805 5776 2839
rect 5724 2796 5776 2805
rect 6000 2796 6052 2848
rect 6644 2796 6696 2848
rect 7104 2796 7156 2848
rect 7564 2839 7616 2848
rect 7564 2805 7573 2839
rect 7573 2805 7607 2839
rect 7607 2805 7616 2839
rect 7564 2796 7616 2805
rect 8024 2839 8076 2848
rect 8024 2805 8033 2839
rect 8033 2805 8067 2839
rect 8067 2805 8076 2839
rect 8024 2796 8076 2805
rect 8484 2796 8536 2848
rect 8668 2839 8720 2848
rect 8668 2805 8677 2839
rect 8677 2805 8711 2839
rect 8711 2805 8720 2839
rect 8668 2796 8720 2805
rect 9404 2796 9456 2848
rect 9588 2796 9640 2848
rect 10324 2839 10376 2848
rect 10324 2805 10333 2839
rect 10333 2805 10367 2839
rect 10367 2805 10376 2839
rect 10324 2796 10376 2805
rect 10784 2839 10836 2848
rect 10784 2805 10793 2839
rect 10793 2805 10827 2839
rect 10827 2805 10836 2839
rect 10784 2796 10836 2805
rect 11244 2796 11296 2848
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 14832 2796 14884 2848
rect 15016 2839 15068 2848
rect 15016 2805 15025 2839
rect 15025 2805 15059 2839
rect 15059 2805 15068 2839
rect 15016 2796 15068 2805
rect 15384 2796 15436 2848
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 16948 2796 17000 2805
rect 18144 2796 18196 2848
rect 18604 2796 18656 2848
rect 19064 2796 19116 2848
rect 19616 2796 19668 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 7288 2592 7340 2644
rect 7656 2635 7708 2644
rect 7656 2601 7665 2635
rect 7665 2601 7699 2635
rect 7699 2601 7708 2635
rect 7656 2592 7708 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 14188 2592 14240 2644
rect 14648 2592 14700 2644
rect 14924 2592 14976 2644
rect 16120 2592 16172 2644
rect 20536 2592 20588 2644
rect 8300 2524 8352 2576
rect 9680 2524 9732 2576
rect 10692 2456 10744 2508
rect 2964 2388 3016 2440
rect 3424 2388 3476 2440
rect 4344 2388 4396 2440
rect 4804 2388 4856 2440
rect 5264 2388 5316 2440
rect 5724 2388 5776 2440
rect 6000 2388 6052 2440
rect 6644 2388 6696 2440
rect 7104 2388 7156 2440
rect 7564 2388 7616 2440
rect 8024 2388 8076 2440
rect 8484 2388 8536 2440
rect 9404 2388 9456 2440
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 10324 2388 10376 2440
rect 10784 2388 10836 2440
rect 11244 2388 11296 2440
rect 13728 2524 13780 2576
rect 14004 2524 14056 2576
rect 15016 2456 15068 2508
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 14188 2388 14240 2440
rect 2044 2252 2096 2304
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 3056 2252 3108 2304
rect 3516 2252 3568 2304
rect 4620 2295 4672 2304
rect 4620 2261 4629 2295
rect 4629 2261 4663 2295
rect 4663 2261 4672 2295
rect 4620 2252 4672 2261
rect 5540 2295 5592 2304
rect 5540 2261 5549 2295
rect 5549 2261 5583 2295
rect 5583 2261 5592 2295
rect 5540 2252 5592 2261
rect 14280 2320 14332 2372
rect 15200 2388 15252 2440
rect 17132 2524 17184 2576
rect 17224 2524 17276 2576
rect 16304 2456 16356 2508
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16856 2388 16908 2440
rect 20076 2456 20128 2508
rect 20352 2456 20404 2508
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18512 2388 18564 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 16028 2320 16080 2372
rect 16304 2320 16356 2372
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 10692 2295 10744 2304
rect 10692 2261 10701 2295
rect 10701 2261 10735 2295
rect 10735 2261 10744 2295
rect 10692 2252 10744 2261
rect 11060 2252 11112 2304
rect 11336 2252 11388 2304
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 12164 2252 12216 2304
rect 12624 2252 12676 2304
rect 13084 2252 13136 2304
rect 13544 2252 13596 2304
rect 14464 2252 14516 2304
rect 15844 2252 15896 2304
rect 17592 2320 17644 2372
rect 17684 2252 17736 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 2320 2048 2372 2100
rect 10692 2048 10744 2100
rect 19524 2048 19576 2100
rect 3056 1980 3108 2032
rect 11060 1980 11112 2032
rect 13820 1980 13872 2032
rect 20260 1980 20312 2032
rect 4620 1912 4672 1964
rect 17960 1912 18012 1964
rect 3516 1844 3568 1896
rect 12348 1844 12400 1896
rect 15108 1844 15160 1896
rect 19248 1844 19300 1896
rect 5540 1776 5592 1828
rect 15936 1776 15988 1828
rect 10232 1708 10284 1760
rect 18052 1708 18104 1760
rect 15568 1640 15620 1692
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 5736 20466 5764 22200
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 7104 20528 7156 20534
rect 17236 20482 17264 22200
rect 20074 21448 20130 21457
rect 20074 21383 20130 21392
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18064 20505 18092 20538
rect 7104 20470 7156 20476
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 1492 11552 1544 11558
rect 1490 11520 1492 11529
rect 1544 11520 1546 11529
rect 1490 11455 1546 11464
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2516 2854 2544 2994
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2056 800 2084 2246
rect 2332 2106 2360 2246
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2516 800 2544 2790
rect 2976 2446 3004 3334
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3896 2854 3924 2994
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3436 2446 3464 2790
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 2976 800 3004 2382
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 2038 3096 2246
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 3436 800 3464 2382
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 1902 3556 2246
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3896 800 3924 2790
rect 4356 2446 4384 3334
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4816 2446 4844 2790
rect 5092 2650 5120 8774
rect 6012 4622 6040 20198
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 7116 19514 7144 20470
rect 17144 20466 17264 20482
rect 18050 20496 18106 20505
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 17132 20460 17264 20466
rect 17184 20454 17264 20460
rect 17316 20460 17368 20466
rect 17132 20402 17184 20408
rect 17316 20402 17368 20408
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17592 20460 17644 20466
rect 20088 20466 20116 21383
rect 20626 21040 20682 21049
rect 20626 20975 20682 20984
rect 20640 20466 20668 20975
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 18050 20431 18106 20440
rect 18144 20460 18196 20466
rect 17592 20402 17644 20408
rect 18144 20402 18196 20408
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8220 19854 8248 20334
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19514 7788 19654
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 7852 12238 7880 19314
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8036 18970 8064 19246
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8404 18766 8432 19110
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18358 8432 18566
rect 8588 18426 8616 20402
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 9140 20058 9168 20402
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9232 20058 9260 20198
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8680 16454 8708 19654
rect 8852 19440 8904 19446
rect 8850 19408 8852 19417
rect 8904 19408 8906 19417
rect 9416 19378 9444 19858
rect 9508 19514 9536 20334
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 9600 19922 9628 20198
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19514 10548 19654
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10888 19446 10916 20198
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 9864 19440 9916 19446
rect 9864 19382 9916 19388
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10876 19440 10928 19446
rect 11060 19440 11112 19446
rect 10876 19382 10928 19388
rect 10980 19388 11060 19394
rect 10980 19382 11112 19388
rect 8850 19343 8906 19352
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9876 19242 9904 19382
rect 10796 19258 10824 19382
rect 10980 19366 11100 19382
rect 10980 19258 11008 19366
rect 11164 19310 11192 19790
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 9864 19236 9916 19242
rect 10796 19230 11008 19258
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 9864 19178 9916 19184
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18426 9260 18566
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9508 18222 9536 18634
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5276 2446 5304 2790
rect 5736 2446 5764 2790
rect 6012 2446 6040 2790
rect 6656 2446 6684 2790
rect 7116 2446 7144 2790
rect 7300 2650 7328 11018
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4282 7512 4422
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7576 2446 7604 2790
rect 7668 2650 7696 8774
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8036 2446 8064 2790
rect 8128 2650 8156 9930
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8312 2582 8340 13874
rect 8496 3194 8524 16390
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 9324 11898 9352 18158
rect 9876 16658 9904 19178
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10520 16794 10548 19110
rect 11164 18766 11192 19246
rect 11256 19174 11284 19722
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11716 18970 11744 20402
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 20058 13124 20198
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13096 19854 13124 19994
rect 13188 19922 13216 20266
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 15120 20058 15148 20198
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 15304 19854 15332 20402
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 16856 19848 16908 19854
rect 16908 19796 16988 19802
rect 16856 19790 16988 19796
rect 16868 19774 16988 19790
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11164 18426 11192 18702
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9416 14006 9444 16594
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15366 9628 16050
rect 10980 15910 11008 16390
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9600 13802 9628 15302
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9876 12306 9904 15846
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10060 12306 10088 14010
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13394 11192 13670
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11256 12306 11284 18906
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11900 18426 11928 18838
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 17338 11744 18362
rect 11900 17678 11928 18362
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11716 16794 11744 17274
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11808 16590 11836 17478
rect 11796 16584 11848 16590
rect 11992 16574 12020 19450
rect 12162 19408 12218 19417
rect 12162 19343 12218 19352
rect 11796 16526 11848 16532
rect 11900 16546 12020 16574
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11716 13258 11744 14214
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8574 4584 8630 4593
rect 8574 4519 8630 4528
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8496 2446 8524 2790
rect 8588 2650 8616 4519
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 9232 3194 9260 8502
rect 9770 6352 9826 6361
rect 9770 6287 9826 6296
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8680 2854 8708 2994
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 4356 800 4384 2382
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4632 1970 4660 2246
rect 4620 1964 4672 1970
rect 4620 1906 4672 1912
rect 4816 800 4844 2382
rect 5276 800 5304 2382
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5552 1834 5580 2246
rect 5540 1828 5592 1834
rect 5540 1770 5592 1776
rect 5736 800 5764 2382
rect 6012 1714 6040 2382
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6012 1686 6224 1714
rect 6196 800 6224 1686
rect 6656 800 6684 2382
rect 7116 800 7144 2382
rect 7576 800 7604 2382
rect 8036 800 8064 2382
rect 8496 800 8524 2382
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8680 762 8708 2790
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9416 2446 9444 2790
rect 9600 2446 9628 2790
rect 9692 2582 9720 5306
rect 9784 2650 9812 6287
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 10336 2446 10364 2790
rect 10704 2514 10732 6122
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10796 2446 10824 2790
rect 11164 2650 11192 10134
rect 11256 2938 11284 12038
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11716 11218 11744 13194
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11808 9654 11836 16526
rect 11900 12442 11928 16546
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 12084 14822 12112 15370
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13870 12020 14350
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12084 12782 12112 14758
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 12176 9450 12204 19343
rect 12636 18698 12664 19654
rect 14936 19514 14964 19654
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 16408 19446 16436 19654
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18766 13860 19110
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11256 2910 11376 2938
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2446 11284 2790
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 8864 870 8984 898
rect 8864 762 8892 870
rect 8956 800 8984 870
rect 9416 800 9444 2382
rect 9600 1714 9628 2382
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 1766 10272 2246
rect 10232 1760 10284 1766
rect 9600 1686 9904 1714
rect 10232 1702 10284 1708
rect 9876 800 9904 1686
rect 10336 800 10364 2382
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10704 2106 10732 2246
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10796 800 10824 2382
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 2038 11100 2246
rect 11060 2032 11112 2038
rect 11060 1974 11112 1980
rect 11256 800 11284 2382
rect 11348 2310 11376 2910
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11716 800 11744 2246
rect 12176 800 12204 2246
rect 12360 1902 12388 11698
rect 12636 11694 12664 18634
rect 15948 18630 15976 19246
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16316 18970 16344 19110
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13188 14804 13216 18226
rect 13280 18086 13308 18566
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13280 17542 13308 18022
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17066 13308 17478
rect 15580 17202 15608 17750
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15856 17270 15884 17478
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13280 16658 13308 17002
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13280 15910 13308 16594
rect 13740 16454 13768 17138
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14568 16522 14596 16934
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13280 15366 13308 15846
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 14958 13308 15302
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13636 14816 13688 14822
rect 13188 14776 13308 14804
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 13190 12848 13874
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 11694 12848 13126
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12452 11286 12480 11630
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12544 2922 12572 9522
rect 12912 9518 12940 14214
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12102 13216 12582
rect 13280 12306 13308 14776
rect 13636 14758 13688 14764
rect 13648 14414 13676 14758
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13648 13734 13676 14350
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13326 13676 13670
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13740 12374 13768 16390
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14074 13860 14962
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 13188 6186 13216 12038
rect 13648 11830 13676 12310
rect 13832 12306 13860 14010
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 14568 13394 14596 16458
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 15026 14872 15302
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14844 14618 14872 14962
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13542 11248 13598 11257
rect 13542 11183 13598 11192
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13358 4040 13414 4049
rect 13358 3975 13414 3984
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 13004 2446 13032 3606
rect 13266 3496 13322 3505
rect 13266 3431 13268 3440
rect 13320 3431 13322 3440
rect 13268 3402 13320 3408
rect 13372 2854 13400 3975
rect 13556 3534 13584 11183
rect 13832 9674 13860 12106
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13740 9646 13860 9674
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13740 2582 13768 9646
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14554 8392 14610 8401
rect 14554 8327 14610 8336
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13924 3058 13952 3402
rect 14292 3074 14320 5578
rect 14384 3534 14412 5782
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14200 3046 14320 3074
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 12636 800 12664 2246
rect 13096 800 13124 2246
rect 13556 800 13584 2246
rect 13832 2038 13860 2926
rect 14200 2922 14228 3046
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14476 2774 14504 4762
rect 14568 3534 14596 8327
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 3097 14596 3334
rect 14554 3088 14610 3097
rect 14554 3023 14610 3032
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14292 2746 14504 2774
rect 14660 2774 14688 5850
rect 14752 4146 14780 12650
rect 15028 12442 15056 12718
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 11354 14872 11630
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10266 15056 10542
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15212 10062 15240 12038
rect 15304 11898 15332 12718
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 10810 15332 10950
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9654 15240 9862
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 8838 15056 9386
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3738 14780 3878
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3058 14780 3470
rect 14844 3466 14872 6054
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15120 4214 15148 4558
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14936 3058 14964 3878
rect 15028 3534 15056 3878
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14830 2952 14886 2961
rect 14830 2887 14886 2896
rect 14844 2854 14872 2887
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14660 2746 14780 2774
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 13820 2032 13872 2038
rect 13820 1974 13872 1980
rect 14016 800 14044 2518
rect 14200 2446 14228 2586
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14292 2378 14320 2746
rect 14648 2644 14700 2650
rect 14752 2632 14780 2746
rect 14700 2604 14780 2632
rect 14924 2644 14976 2650
rect 14648 2586 14700 2592
rect 14924 2586 14976 2592
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 800 14504 2246
rect 14936 800 14964 2586
rect 15028 2514 15056 2790
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15120 1902 15148 4150
rect 15212 2446 15240 4694
rect 15304 3534 15332 7414
rect 15396 4146 15424 12038
rect 15488 11898 15516 12174
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15580 10130 15608 17138
rect 15856 16590 15884 17206
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15856 15570 15884 16186
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15948 15450 15976 18566
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16960 18358 16988 19774
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16776 18170 16804 18226
rect 16316 17542 16344 18158
rect 16776 18142 16988 18170
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16212 16516 16264 16522
rect 16212 16458 16264 16464
rect 15856 15422 15976 15450
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 10810 15700 11698
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15488 8294 15516 9998
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 9178 15608 9454
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15764 7546 15792 13942
rect 15856 12306 15884 15422
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 12866 15976 14350
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16224 13818 16252 16458
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16960 15910 16988 18142
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16316 15162 16344 15506
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16316 14414 16344 15098
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16304 14408 16356 14414
rect 16684 14385 16712 14758
rect 16304 14350 16356 14356
rect 16670 14376 16726 14385
rect 16316 13938 16344 14350
rect 16670 14311 16726 14320
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16960 14074 16988 14282
rect 17144 14226 17172 18634
rect 17328 18426 17356 20402
rect 17512 19922 17540 20402
rect 17604 19990 17632 20402
rect 17958 20360 18014 20369
rect 17958 20295 17960 20304
rect 18012 20295 18014 20304
rect 17960 20266 18012 20272
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 18834 17632 19654
rect 18064 19378 18092 20198
rect 18156 19514 18184 20402
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18248 19825 18276 20198
rect 18234 19816 18290 19825
rect 18234 19751 18290 19760
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17224 14340 17276 14346
rect 17328 14328 17356 17002
rect 17512 16454 17540 18226
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17276 14300 17356 14328
rect 17224 14282 17276 14288
rect 17052 14198 17172 14226
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16040 13326 16068 13806
rect 16224 13790 16344 13818
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 12986 16160 13262
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15948 12838 16160 12866
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16040 11558 16068 12038
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15856 9110 15884 11154
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10198 15976 10406
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15580 3126 15608 7278
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15672 4146 15700 6122
rect 15764 5778 15792 7482
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15948 4690 15976 5170
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16040 4570 16068 11494
rect 16132 9042 16160 12838
rect 16224 12442 16252 13126
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16316 9042 16344 13790
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12238 16436 13126
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12374 16988 12582
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 17052 12306 17080 14198
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16946 11792 17002 11801
rect 16946 11727 17002 11736
rect 16960 11626 16988 11727
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16868 11286 16896 11494
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16960 10062 16988 10950
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 8430 16344 8978
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15948 4542 16068 4570
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15856 3194 15884 3878
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15396 800 15424 2790
rect 15580 1698 15608 2926
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15764 2446 15792 2858
rect 15948 2774 15976 4542
rect 16132 4146 16160 8298
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16316 5370 16344 7754
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4214 16344 4422
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16040 3126 16068 3470
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 15856 2746 15976 2774
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15856 2394 15884 2746
rect 15856 2366 15976 2394
rect 16040 2378 16068 2790
rect 16132 2650 16160 2994
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16316 2514 16344 3878
rect 16408 3534 16436 4966
rect 16960 4622 16988 9862
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 17052 4468 17080 11494
rect 17144 10606 17172 13670
rect 17236 13190 17264 13942
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17236 10198 17264 13126
rect 17328 10810 17356 14300
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17144 8498 17172 8774
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16960 4440 17080 4468
rect 17132 4480 17184 4486
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16960 4196 16988 4440
rect 17132 4422 17184 4428
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 16486 4176 16542 4185
rect 16868 4168 16988 4196
rect 16486 4111 16542 4120
rect 16764 4140 16816 4146
rect 16500 3738 16528 4111
rect 16764 4082 16816 4088
rect 16776 4010 16804 4082
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16868 3534 16896 4168
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3058 16436 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16960 3074 16988 3538
rect 17052 3534 17080 4218
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16868 3046 16988 3074
rect 17144 3058 17172 4422
rect 17236 4026 17264 9930
rect 17328 9178 17356 10610
rect 17420 10130 17448 15846
rect 17512 13734 17540 16390
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17604 12782 17632 18770
rect 17972 18630 18000 19110
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18154 18000 18566
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 17678 18000 18090
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17972 17270 18000 17614
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 14074 17724 16934
rect 17972 16590 18000 17206
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17512 12102 17540 12310
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17512 11626 17540 12038
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17512 10146 17540 11562
rect 17604 11506 17632 11834
rect 17696 11694 17724 14010
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17604 11478 17816 11506
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 10266 17632 11086
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17408 10124 17460 10130
rect 17512 10118 17632 10146
rect 17408 10066 17460 10072
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9722 17540 9998
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8566 17540 8774
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17328 5658 17356 6802
rect 17512 6798 17540 7142
rect 17604 6866 17632 10118
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17420 5778 17448 6598
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17328 5630 17448 5658
rect 17314 5400 17370 5409
rect 17314 5335 17370 5344
rect 17328 5302 17356 5335
rect 17316 5296 17368 5302
rect 17316 5238 17368 5244
rect 17328 5166 17356 5238
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17314 4176 17370 4185
rect 17314 4111 17316 4120
rect 17368 4111 17370 4120
rect 17316 4082 17368 4088
rect 17236 3998 17356 4026
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17132 3052 17184 3058
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 16868 2446 16896 3046
rect 17132 2994 17184 3000
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15568 1692 15620 1698
rect 15568 1634 15620 1640
rect 15856 800 15884 2246
rect 15948 1834 15976 2366
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 15936 1828 15988 1834
rect 15936 1770 15988 1776
rect 16316 800 16344 2314
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 1442 16988 2790
rect 17236 2666 17264 3878
rect 17328 3738 17356 3998
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17420 2990 17448 5630
rect 17512 4486 17540 6258
rect 17604 5370 17632 6598
rect 17696 5710 17724 11290
rect 17788 9761 17816 11478
rect 17880 11354 17908 16458
rect 18064 16402 18092 18022
rect 18524 17202 18552 19450
rect 18800 19417 18828 20198
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 21376 19922 21404 20334
rect 22468 20324 22520 20330
rect 22468 20266 22520 20272
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 18786 19408 18842 19417
rect 18786 19343 18842 19352
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16794 18552 17138
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 17972 16374 18092 16402
rect 17972 16114 18000 16374
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 16017 18000 16050
rect 18052 16040 18104 16046
rect 17958 16008 18014 16017
rect 18052 15982 18104 15988
rect 17958 15943 18014 15952
rect 18064 15570 18092 15982
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 18064 15026 18092 15506
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18248 14822 18276 15370
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17972 12238 18000 13194
rect 18064 12434 18092 14554
rect 18156 13258 18184 14758
rect 18340 14278 18368 15098
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18156 13138 18184 13194
rect 18156 13110 18276 13138
rect 18064 12406 18184 12434
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 18064 11218 18092 11698
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17868 10736 17920 10742
rect 17972 10713 18000 11018
rect 17868 10678 17920 10684
rect 17958 10704 18014 10713
rect 17774 9752 17830 9761
rect 17774 9687 17830 9696
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17788 8090 17816 9522
rect 17880 9450 17908 10678
rect 17958 10639 18014 10648
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17866 9344 17922 9353
rect 17866 9279 17922 9288
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17880 7698 17908 9279
rect 17972 8634 18000 10474
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 7993 18000 8434
rect 17958 7984 18014 7993
rect 17958 7919 18014 7928
rect 17788 7670 17908 7698
rect 17788 6662 17816 7670
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17880 7449 17908 7482
rect 17866 7440 17922 7449
rect 17866 7375 17922 7384
rect 18064 7342 18092 8774
rect 18156 7954 18184 12406
rect 18248 10146 18276 13110
rect 18340 10418 18368 14214
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18432 13977 18460 14010
rect 18418 13968 18474 13977
rect 18524 13938 18552 14350
rect 18418 13903 18474 13912
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18524 13394 18552 13874
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18616 12434 18644 17614
rect 18708 12986 18736 18702
rect 18892 17882 18920 19450
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19628 19009 19656 19654
rect 19614 19000 19670 19009
rect 19614 18935 19670 18944
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19168 18290 19196 18566
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 17134 19288 17614
rect 19248 17128 19300 17134
rect 18970 17096 19026 17105
rect 19248 17070 19300 17076
rect 18970 17031 18972 17040
rect 19024 17031 19026 17040
rect 18972 17002 19024 17008
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18524 12406 18644 12434
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11354 18460 12038
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18524 10810 18552 12406
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18616 10606 18644 12038
rect 18800 11694 18828 16730
rect 19248 16584 19300 16590
rect 19154 16552 19210 16561
rect 19248 16526 19300 16532
rect 19154 16487 19210 16496
rect 19168 16250 19196 16487
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19260 16046 19288 16526
rect 19536 16522 19564 18226
rect 19614 18184 19670 18193
rect 19614 18119 19616 18128
rect 19668 18119 19670 18128
rect 19616 18090 19668 18096
rect 19720 17542 19748 19722
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 17610 19932 18566
rect 20272 18290 20300 19110
rect 20640 18737 20668 19110
rect 20626 18728 20682 18737
rect 20352 18692 20404 18698
rect 20626 18663 20682 18672
rect 20352 18634 20404 18640
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20272 18170 20300 18226
rect 20180 18142 20300 18170
rect 19892 17604 19944 17610
rect 19892 17546 19944 17552
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19246 15464 19302 15473
rect 19246 15399 19302 15408
rect 19260 15366 19288 15399
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19522 14920 19578 14929
rect 19522 14855 19578 14864
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18340 10390 18644 10418
rect 18248 10118 18460 10146
rect 18236 10056 18288 10062
rect 18234 10024 18236 10033
rect 18288 10024 18290 10033
rect 18234 9959 18290 9968
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18248 9722 18276 9862
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 8498 18276 9522
rect 18340 9178 18368 9862
rect 18432 9518 18460 10118
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18432 9042 18460 9454
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 6866 18092 7142
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6322 17816 6598
rect 18156 6458 18184 7686
rect 18340 7562 18368 8910
rect 18510 8664 18566 8673
rect 18510 8599 18566 8608
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18248 7534 18368 7562
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17972 6225 18000 6258
rect 17958 6216 18014 6225
rect 17958 6151 18014 6160
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17696 2774 17724 4762
rect 17788 4622 17816 6054
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17880 4729 17908 5782
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17972 5545 18000 5578
rect 17958 5536 18014 5545
rect 17958 5471 18014 5480
rect 18064 5137 18092 6326
rect 18248 5710 18276 7534
rect 18432 7478 18460 7686
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18340 7313 18368 7346
rect 18326 7304 18382 7313
rect 18326 7239 18382 7248
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18340 6361 18368 6734
rect 18326 6352 18382 6361
rect 18524 6322 18552 8599
rect 18616 6934 18644 10390
rect 18708 10266 18736 10610
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18694 8392 18750 8401
rect 18694 8327 18696 8336
rect 18748 8327 18750 8336
rect 18696 8298 18748 8304
rect 18800 8090 18828 8434
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18326 6287 18382 6296
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18050 5128 18106 5137
rect 18050 5063 18106 5072
rect 17866 4720 17922 4729
rect 17866 4655 17922 4664
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 4185 18000 4490
rect 17958 4176 18014 4185
rect 17958 4111 18014 4120
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17144 2638 17264 2666
rect 17604 2746 17724 2774
rect 17144 2582 17172 2638
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 16776 1414 16988 1442
rect 16776 800 16804 1414
rect 17236 800 17264 2518
rect 17604 2378 17632 2746
rect 17788 2446 17816 3878
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 800 17724 2246
rect 17972 1970 18000 3334
rect 17960 1964 18012 1970
rect 17960 1906 18012 1912
rect 18064 1766 18092 4014
rect 18156 3058 18184 5510
rect 18524 5166 18552 6258
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 5914 18644 6190
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18248 4282 18276 5102
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18234 3632 18290 3641
rect 18234 3567 18236 3576
rect 18288 3567 18290 3576
rect 18236 3538 18288 3544
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 18156 800 18184 2790
rect 18524 2446 18552 4966
rect 18708 4758 18736 7958
rect 18892 7478 18920 13942
rect 18984 13433 19012 14758
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19536 14618 19564 14855
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19720 14498 19748 17138
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19812 14822 19840 16050
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19628 14470 19748 14498
rect 19628 14074 19656 14470
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 18970 13424 19026 13433
rect 18970 13359 19026 13368
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18984 12442 19012 12854
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 19076 11898 19104 12650
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19720 12442 19748 14350
rect 19708 12436 19760 12442
rect 19812 12434 19840 14758
rect 19904 12782 19932 17546
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 14006 20024 15302
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13394 20024 13670
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 20088 13326 20116 16390
rect 20076 13320 20128 13326
rect 19982 13288 20038 13297
rect 20076 13262 20128 13268
rect 19982 13223 20038 13232
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19812 12406 19932 12434
rect 19708 12378 19760 12384
rect 19154 12336 19210 12345
rect 19154 12271 19210 12280
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19168 11778 19196 12271
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19536 11898 19564 12106
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19076 11750 19196 11778
rect 19616 11756 19668 11762
rect 19076 11218 19104 11750
rect 19616 11698 19668 11704
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19536 11354 19564 11494
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10810 19380 11086
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19628 10554 19656 11698
rect 19536 10526 19656 10554
rect 19536 10470 19564 10526
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 18972 8968 19024 8974
rect 18970 8936 18972 8945
rect 19024 8936 19026 8945
rect 19026 8894 19104 8922
rect 18970 8871 19026 8880
rect 18970 8392 19026 8401
rect 18970 8327 19026 8336
rect 18984 7886 19012 8327
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19076 7478 19104 8894
rect 19260 8498 19288 9007
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19352 8634 19380 8774
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19536 7546 19564 9522
rect 19628 8838 19656 9590
rect 19720 9058 19748 11834
rect 19812 11354 19840 12038
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19904 10826 19932 12406
rect 19996 11694 20024 13223
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19996 11257 20024 11290
rect 19982 11248 20038 11257
rect 19982 11183 20038 11192
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19812 10798 19932 10826
rect 19812 9194 19840 10798
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19904 9722 19932 10610
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19812 9166 19932 9194
rect 19996 9178 20024 11086
rect 20088 10198 20116 12174
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 20180 10146 20208 18142
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 12306 20300 17478
rect 20364 13433 20392 18634
rect 20720 18624 20772 18630
rect 20640 18572 20720 18578
rect 20640 18566 20772 18572
rect 20640 18550 20760 18566
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20350 13424 20406 13433
rect 20350 13359 20406 13368
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20258 12200 20314 12209
rect 20258 12135 20314 12144
rect 20272 11150 20300 12135
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20364 10826 20392 13194
rect 20456 11626 20484 17206
rect 20548 16153 20576 17478
rect 20640 17241 20668 18550
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20626 17232 20682 17241
rect 20626 17167 20682 17176
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20534 16144 20590 16153
rect 20534 16079 20590 16088
rect 20640 15745 20668 17002
rect 20732 16998 20760 17818
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20824 16522 20852 19654
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 17785 21312 19110
rect 21560 18086 21588 19722
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21270 17776 21326 17785
rect 21270 17711 21326 17720
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20626 15736 20682 15745
rect 20626 15671 20682 15680
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20640 15094 20668 15438
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20640 14414 20668 15030
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20732 14226 20760 16118
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20824 14278 20852 14962
rect 21008 14346 21036 15846
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20640 14198 20760 14226
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20364 10798 20484 10826
rect 20548 10810 20576 13874
rect 20640 13870 20668 14198
rect 21008 14090 21036 14282
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20824 14062 21036 14090
rect 20732 13977 20760 14010
rect 20718 13968 20774 13977
rect 20718 13903 20774 13912
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20180 10118 20300 10146
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20180 9722 20208 9930
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19720 9030 19840 9058
rect 19904 9042 19932 9166
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19628 8514 19656 8774
rect 19720 8634 19748 8910
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19628 8486 19748 8514
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18800 4010 18828 7346
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18892 4010 18920 7278
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 18972 6792 19024 6798
rect 18970 6760 18972 6769
rect 19024 6760 19026 6769
rect 18970 6695 19026 6704
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 18984 5234 19012 6598
rect 19260 6458 19288 6598
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19444 6202 19472 6938
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19536 6730 19564 6802
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19444 6174 19564 6202
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19536 5794 19564 6174
rect 19444 5766 19564 5794
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19260 5302 19288 5510
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19444 5098 19472 5766
rect 19522 5672 19578 5681
rect 19522 5607 19578 5616
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19444 4554 19472 4762
rect 19536 4690 19564 5607
rect 19628 5166 19656 7890
rect 19720 7886 19748 8486
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19720 7449 19748 7482
rect 19706 7440 19762 7449
rect 19706 7375 19762 7384
rect 19720 5370 19748 7375
rect 19812 6866 19840 9030
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 20272 8650 20300 10118
rect 20364 9450 20392 10610
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20088 8622 20300 8650
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19904 7750 19932 8230
rect 20088 7954 20116 8622
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19904 7002 19932 7686
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19812 5658 19840 6802
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19904 5778 19932 6666
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19812 5630 19932 5658
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19616 5160 19668 5166
rect 19668 5108 19748 5114
rect 19616 5102 19748 5108
rect 19628 5086 19748 5102
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19614 4584 19670 4593
rect 19432 4548 19484 4554
rect 19614 4519 19616 4528
rect 19432 4490 19484 4496
rect 19668 4519 19670 4528
rect 19616 4490 19668 4496
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19352 4282 19380 4422
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18604 3528 18656 3534
rect 18602 3496 18604 3505
rect 18656 3496 18658 3505
rect 18602 3431 18658 3440
rect 18786 3496 18842 3505
rect 18786 3431 18788 3440
rect 18840 3431 18842 3440
rect 18788 3402 18840 3408
rect 19076 3194 19104 3878
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19536 3602 19564 4422
rect 19720 3602 19748 5086
rect 19812 4554 19840 5510
rect 19904 4826 19932 5630
rect 19996 5234 20024 6870
rect 20088 6866 20116 7686
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20180 6662 20208 8366
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20088 5574 20116 6598
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 19800 4548 19852 4554
rect 19800 4490 19852 4496
rect 19996 4298 20024 5034
rect 19904 4270 20024 4298
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19812 3602 19840 4150
rect 19904 3618 19932 4270
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19996 4049 20024 4082
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 20088 3738 20116 5306
rect 20272 5098 20300 8502
rect 20364 8090 20392 8774
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20350 7440 20406 7449
rect 20350 7375 20406 7384
rect 20364 6322 20392 7375
rect 20456 6338 20484 10798
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20640 10538 20668 12786
rect 20732 11830 20760 13126
rect 20824 12714 20852 14062
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20916 12434 20944 12786
rect 20824 12406 20944 12434
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20824 10810 20852 12406
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20824 10266 20852 10610
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20548 6458 20576 9522
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20640 9178 20668 9454
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20640 7410 20668 8842
rect 20732 8634 20760 9862
rect 20916 9518 20944 12310
rect 21008 10810 21036 13874
rect 21100 12986 21128 17138
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 21100 12374 21128 12650
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20640 6934 20668 7346
rect 20732 7274 20760 7890
rect 20824 7546 20852 8774
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20352 6316 20404 6322
rect 20456 6310 20576 6338
rect 20352 6258 20404 6264
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20364 4826 20392 6258
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20456 5914 20484 6190
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20180 4146 20208 4762
rect 20456 4486 20484 5578
rect 20548 4690 20576 6310
rect 20640 5370 20668 6598
rect 20732 5778 20760 7210
rect 20810 6488 20866 6497
rect 20810 6423 20866 6432
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20824 5710 20852 6423
rect 20916 6254 20944 8978
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20260 4480 20312 4486
rect 20444 4480 20496 4486
rect 20260 4422 20312 4428
rect 20364 4428 20444 4434
rect 20364 4422 20496 4428
rect 20272 4282 20300 4422
rect 20364 4406 20484 4422
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19800 3596 19852 3602
rect 19904 3590 20116 3618
rect 19800 3538 19852 3544
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19338 3088 19394 3097
rect 19338 3023 19340 3032
rect 19392 3023 19394 3032
rect 19340 2994 19392 3000
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18616 800 18644 2790
rect 19076 800 19104 2790
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19536 2106 19564 3402
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19904 2961 19932 2994
rect 19890 2952 19946 2961
rect 19890 2887 19946 2896
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19524 2100 19576 2106
rect 19524 2042 19576 2048
rect 19248 1896 19300 1902
rect 19248 1838 19300 1844
rect 19260 1465 19288 1838
rect 19246 1456 19302 1465
rect 19628 1442 19656 2790
rect 19246 1391 19302 1400
rect 19536 1414 19656 1442
rect 19536 800 19564 1414
rect 19996 800 20024 3334
rect 20088 2514 20116 3590
rect 20180 3398 20208 3946
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20364 2514 20392 4406
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 3913 20576 4014
rect 20534 3904 20590 3913
rect 20534 3839 20590 3848
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20548 3097 20576 3470
rect 20534 3088 20590 3097
rect 20640 3058 20668 5170
rect 20732 3602 20760 5510
rect 20824 4214 20852 5510
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20916 3738 20944 5102
rect 21008 4758 21036 9862
rect 21100 9178 21128 12174
rect 21192 11354 21220 17614
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 14521 21312 16390
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21270 14512 21326 14521
rect 21270 14447 21326 14456
rect 21272 13728 21324 13734
rect 21270 13696 21272 13705
rect 21324 13696 21326 13705
rect 21270 13631 21326 13640
rect 21376 13530 21404 15302
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21468 14006 21496 14894
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21270 13288 21326 13297
rect 21270 13223 21326 13232
rect 21284 12986 21312 13223
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21270 12880 21326 12889
rect 21270 12815 21326 12824
rect 21284 12442 21312 12815
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21192 8022 21220 9318
rect 21284 8634 21312 11630
rect 21376 11150 21404 12582
rect 21468 11898 21496 13806
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21454 11248 21510 11257
rect 21454 11183 21510 11192
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21468 11082 21496 11183
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21468 10810 21496 11018
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21362 10432 21418 10441
rect 21362 10367 21418 10376
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21376 8498 21404 10367
rect 21454 9616 21510 9625
rect 21454 9551 21510 9560
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21100 5166 21128 6802
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20534 3023 20590 3032
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20272 2038 20300 2382
rect 20260 2032 20312 2038
rect 20260 1974 20312 1980
rect 20272 1873 20300 1974
rect 20258 1864 20314 1873
rect 20258 1799 20314 1808
rect 20456 800 20484 2858
rect 20548 2689 20576 2926
rect 20534 2680 20590 2689
rect 20534 2615 20536 2624
rect 20588 2615 20590 2624
rect 20536 2586 20588 2592
rect 20548 2555 20576 2586
rect 20536 2440 20588 2446
rect 20534 2408 20536 2417
rect 20588 2408 20590 2417
rect 20534 2343 20590 2352
rect 20916 800 20944 3538
rect 21192 3194 21220 7142
rect 21284 5574 21312 8298
rect 21468 7410 21496 9551
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21560 6866 21588 18022
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21652 11286 21680 15642
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21730 11656 21786 11665
rect 21730 11591 21786 11600
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21744 11098 21772 11591
rect 21652 11070 21772 11098
rect 21652 9586 21680 11070
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 22112 8430 22140 16458
rect 22204 11558 22232 16526
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22296 7954 22324 13942
rect 22388 10470 22416 18702
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22480 7886 22508 20266
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21362 6760 21418 6769
rect 21362 6695 21364 6704
rect 21416 6695 21418 6704
rect 21364 6666 21416 6672
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 22572 3942 22600 13466
rect 22664 6662 22692 14214
rect 22756 10130 22784 16934
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 8680 734 8892 762
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
<< via2 >>
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 20074 21392 20130 21448
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 1490 11500 1492 11520
rect 1492 11500 1544 11520
rect 1544 11500 1546 11520
rect 1490 11464 1546 11500
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 18050 20440 18106 20496
rect 20626 20984 20682 21040
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8850 19388 8852 19408
rect 8852 19388 8904 19408
rect 8904 19388 8906 19408
rect 8850 19352 8906 19388
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 12162 19352 12218 19408
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8574 4528 8630 4584
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9770 6296 9826 6352
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13542 11192 13598 11248
rect 13358 3984 13414 4040
rect 13266 3460 13322 3496
rect 13266 3440 13268 3460
rect 13268 3440 13320 3460
rect 13320 3440 13322 3460
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14554 8336 14610 8392
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14554 3032 14610 3088
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14830 2896 14886 2952
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16670 14320 16726 14376
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 17958 20324 18014 20360
rect 17958 20304 17960 20324
rect 17960 20304 18012 20324
rect 18012 20304 18014 20324
rect 18234 19760 18290 19816
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16946 11736 17002 11792
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16486 4120 16542 4176
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17314 5344 17370 5400
rect 17314 4140 17370 4176
rect 17314 4120 17316 4140
rect 17316 4120 17368 4140
rect 17368 4120 17370 4140
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 18786 19352 18842 19408
rect 17958 15952 18014 16008
rect 17774 9696 17830 9752
rect 17958 10648 18014 10704
rect 17866 9288 17922 9344
rect 17958 7928 18014 7984
rect 17866 7384 17922 7440
rect 18418 13912 18474 13968
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19614 18944 19670 19000
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 18970 17060 19026 17096
rect 18970 17040 18972 17060
rect 18972 17040 19024 17060
rect 19024 17040 19026 17060
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19154 16496 19210 16552
rect 19614 18148 19670 18184
rect 19614 18128 19616 18148
rect 19616 18128 19668 18148
rect 19668 18128 19670 18148
rect 20626 18672 20682 18728
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19246 15408 19302 15464
rect 19522 14864 19578 14920
rect 18234 10004 18236 10024
rect 18236 10004 18288 10024
rect 18288 10004 18290 10024
rect 18234 9968 18290 10004
rect 18510 8608 18566 8664
rect 17958 6160 18014 6216
rect 17958 5480 18014 5536
rect 18326 7248 18382 7304
rect 18326 6296 18382 6352
rect 18694 8356 18750 8392
rect 18694 8336 18696 8356
rect 18696 8336 18748 8356
rect 18748 8336 18750 8356
rect 18050 5072 18106 5128
rect 17866 4664 17922 4720
rect 17958 4120 18014 4176
rect 18234 3596 18290 3632
rect 18234 3576 18236 3596
rect 18236 3576 18288 3596
rect 18288 3576 18290 3596
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 18970 13368 19026 13424
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19982 13232 20038 13288
rect 19154 12280 19210 12336
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19246 9016 19302 9072
rect 18970 8916 18972 8936
rect 18972 8916 19024 8936
rect 19024 8916 19026 8936
rect 18970 8880 19026 8916
rect 18970 8336 19026 8392
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19982 11192 20038 11248
rect 20350 13368 20406 13424
rect 20258 12144 20314 12200
rect 20626 17176 20682 17232
rect 20534 16088 20590 16144
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21270 17720 21326 17776
rect 20626 15680 20682 15736
rect 20718 13912 20774 13968
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18970 6740 18972 6760
rect 18972 6740 19024 6760
rect 19024 6740 19026 6760
rect 18970 6704 19026 6740
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19522 5616 19578 5672
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19706 7384 19762 7440
rect 19614 4548 19670 4584
rect 19614 4528 19616 4548
rect 19616 4528 19668 4548
rect 19668 4528 19670 4548
rect 18602 3476 18604 3496
rect 18604 3476 18656 3496
rect 18656 3476 18658 3496
rect 18602 3440 18658 3476
rect 18786 3460 18842 3496
rect 18786 3440 18788 3460
rect 18788 3440 18840 3460
rect 18840 3440 18842 3460
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19982 3984 20038 4040
rect 20350 7384 20406 7440
rect 20810 6432 20866 6488
rect 19338 3052 19394 3088
rect 19338 3032 19340 3052
rect 19340 3032 19392 3052
rect 19392 3032 19394 3052
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19890 2896 19946 2952
rect 19246 1400 19302 1456
rect 20534 3848 20590 3904
rect 20534 3032 20590 3088
rect 21270 14456 21326 14512
rect 21270 13676 21272 13696
rect 21272 13676 21324 13696
rect 21324 13676 21326 13696
rect 21270 13640 21326 13676
rect 21270 13232 21326 13288
rect 21270 12824 21326 12880
rect 21454 11192 21510 11248
rect 21362 10376 21418 10432
rect 21454 9560 21510 9616
rect 20258 1808 20314 1864
rect 20534 2644 20590 2680
rect 20534 2624 20536 2644
rect 20536 2624 20588 2644
rect 20588 2624 20590 2644
rect 20534 2388 20536 2408
rect 20536 2388 20588 2408
rect 20588 2388 20590 2408
rect 20534 2352 20590 2388
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21730 11600 21786 11656
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21362 6724 21418 6760
rect 21362 6704 21364 6724
rect 21364 6704 21416 6724
rect 21416 6704 21418 6724
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 20069 21450 20135 21453
rect 22200 21450 23000 21480
rect 20069 21448 23000 21450
rect 20069 21392 20074 21448
rect 20130 21392 23000 21448
rect 20069 21390 23000 21392
rect 20069 21387 20135 21390
rect 22200 21360 23000 21390
rect 20621 21042 20687 21045
rect 22200 21042 23000 21072
rect 20621 21040 23000 21042
rect 20621 20984 20626 21040
rect 20682 20984 23000 21040
rect 20621 20982 23000 20984
rect 20621 20979 20687 20982
rect 22200 20952 23000 20982
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 22200 20634 23000 20664
rect 22142 20544 23000 20634
rect 18045 20498 18111 20501
rect 22142 20498 22202 20544
rect 18045 20496 22202 20498
rect 18045 20440 18050 20496
rect 18106 20440 22202 20496
rect 18045 20438 22202 20440
rect 18045 20435 18111 20438
rect 17953 20362 18019 20365
rect 17953 20360 19994 20362
rect 17953 20304 17958 20360
rect 18014 20304 19994 20360
rect 17953 20302 19994 20304
rect 17953 20299 18019 20302
rect 19934 20226 19994 20302
rect 22200 20226 23000 20256
rect 19934 20166 23000 20226
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 22200 20136 23000 20166
rect 19139 20095 19455 20096
rect 18229 19818 18295 19821
rect 22200 19818 23000 19848
rect 18229 19816 23000 19818
rect 18229 19760 18234 19816
rect 18290 19760 23000 19816
rect 18229 19758 23000 19760
rect 18229 19755 18295 19758
rect 22200 19728 23000 19758
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 8845 19410 8911 19413
rect 12157 19410 12223 19413
rect 8845 19408 12223 19410
rect 8845 19352 8850 19408
rect 8906 19352 12162 19408
rect 12218 19352 12223 19408
rect 8845 19350 12223 19352
rect 8845 19347 8911 19350
rect 12157 19347 12223 19350
rect 18781 19410 18847 19413
rect 22200 19410 23000 19440
rect 18781 19408 23000 19410
rect 18781 19352 18786 19408
rect 18842 19352 23000 19408
rect 18781 19350 23000 19352
rect 18781 19347 18847 19350
rect 22200 19320 23000 19350
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 19609 19002 19675 19005
rect 22200 19002 23000 19032
rect 19609 19000 23000 19002
rect 19609 18944 19614 19000
rect 19670 18944 23000 19000
rect 19609 18942 23000 18944
rect 19609 18939 19675 18942
rect 22200 18912 23000 18942
rect 20621 18730 20687 18733
rect 20621 18728 22202 18730
rect 20621 18672 20626 18728
rect 20682 18672 22202 18728
rect 20621 18670 22202 18672
rect 20621 18667 20687 18670
rect 22142 18624 22202 18670
rect 22142 18534 23000 18624
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 19609 18186 19675 18189
rect 22200 18186 23000 18216
rect 19609 18184 23000 18186
rect 19609 18128 19614 18184
rect 19670 18128 23000 18184
rect 19609 18126 23000 18128
rect 19609 18123 19675 18126
rect 22200 18096 23000 18126
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 21265 17778 21331 17781
rect 22200 17778 23000 17808
rect 21265 17776 23000 17778
rect 21265 17720 21270 17776
rect 21326 17720 23000 17776
rect 21265 17718 23000 17720
rect 21265 17715 21331 17718
rect 22200 17688 23000 17718
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 22200 17370 23000 17400
rect 22142 17280 23000 17370
rect 20621 17234 20687 17237
rect 22142 17234 22202 17280
rect 20621 17232 22202 17234
rect 20621 17176 20626 17232
rect 20682 17176 22202 17232
rect 20621 17174 22202 17176
rect 20621 17171 20687 17174
rect 18965 17098 19031 17101
rect 18965 17096 20730 17098
rect 18965 17040 18970 17096
rect 19026 17040 20730 17096
rect 18965 17038 20730 17040
rect 18965 17035 19031 17038
rect 20670 16962 20730 17038
rect 22200 16962 23000 16992
rect 20670 16902 23000 16962
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 19149 16554 19215 16557
rect 22200 16554 23000 16584
rect 19149 16552 23000 16554
rect 19149 16496 19154 16552
rect 19210 16496 23000 16552
rect 19149 16494 23000 16496
rect 19149 16491 19215 16494
rect 22200 16464 23000 16494
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 20529 16146 20595 16149
rect 22200 16146 23000 16176
rect 20529 16144 23000 16146
rect 20529 16088 20534 16144
rect 20590 16088 23000 16144
rect 20529 16086 23000 16088
rect 20529 16083 20595 16086
rect 22200 16056 23000 16086
rect 17953 16010 18019 16013
rect 18270 16010 18276 16012
rect 17953 16008 18276 16010
rect 17953 15952 17958 16008
rect 18014 15952 18276 16008
rect 17953 15950 18276 15952
rect 17953 15947 18019 15950
rect 18270 15948 18276 15950
rect 18340 15948 18346 16012
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 20621 15738 20687 15741
rect 22200 15738 23000 15768
rect 20621 15736 23000 15738
rect 20621 15680 20626 15736
rect 20682 15680 23000 15736
rect 20621 15678 23000 15680
rect 20621 15675 20687 15678
rect 22200 15648 23000 15678
rect 19241 15466 19307 15469
rect 19241 15464 22202 15466
rect 19241 15408 19246 15464
rect 19302 15408 22202 15464
rect 19241 15406 22202 15408
rect 19241 15403 19307 15406
rect 22142 15360 22202 15406
rect 22142 15270 23000 15360
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 19517 14922 19583 14925
rect 22200 14922 23000 14952
rect 19517 14920 23000 14922
rect 19517 14864 19522 14920
rect 19578 14864 23000 14920
rect 19517 14862 23000 14864
rect 19517 14859 19583 14862
rect 22200 14832 23000 14862
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 21265 14514 21331 14517
rect 22200 14514 23000 14544
rect 21265 14512 23000 14514
rect 21265 14456 21270 14512
rect 21326 14456 23000 14512
rect 21265 14454 23000 14456
rect 21265 14451 21331 14454
rect 22200 14424 23000 14454
rect 16665 14378 16731 14381
rect 17350 14378 17356 14380
rect 16665 14376 17356 14378
rect 16665 14320 16670 14376
rect 16726 14320 17356 14376
rect 16665 14318 17356 14320
rect 16665 14315 16731 14318
rect 17350 14316 17356 14318
rect 17420 14316 17426 14380
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 22200 14106 23000 14136
rect 22142 14016 23000 14106
rect 18413 13972 18479 13973
rect 18413 13968 18460 13972
rect 18524 13970 18530 13972
rect 20713 13970 20779 13973
rect 22142 13970 22202 14016
rect 18413 13912 18418 13968
rect 18413 13908 18460 13912
rect 18524 13910 18570 13970
rect 20713 13968 22202 13970
rect 20713 13912 20718 13968
rect 20774 13912 22202 13968
rect 20713 13910 22202 13912
rect 18524 13908 18530 13910
rect 18413 13907 18479 13908
rect 20713 13907 20779 13910
rect 21265 13698 21331 13701
rect 22200 13698 23000 13728
rect 21265 13696 23000 13698
rect 21265 13640 21270 13696
rect 21326 13640 23000 13696
rect 21265 13638 23000 13640
rect 21265 13635 21331 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22200 13608 23000 13638
rect 19139 13567 19455 13568
rect 18965 13428 19031 13429
rect 18965 13426 19012 13428
rect 18920 13424 19012 13426
rect 18920 13368 18970 13424
rect 18920 13366 19012 13368
rect 18965 13364 19012 13366
rect 19076 13364 19082 13428
rect 20345 13426 20411 13429
rect 20302 13424 20411 13426
rect 20302 13368 20350 13424
rect 20406 13368 20411 13424
rect 18965 13363 19031 13364
rect 20302 13363 20411 13368
rect 19977 13290 20043 13293
rect 20302 13290 20362 13363
rect 19977 13288 20362 13290
rect 19977 13232 19982 13288
rect 20038 13232 20362 13288
rect 19977 13230 20362 13232
rect 21265 13290 21331 13293
rect 22200 13290 23000 13320
rect 21265 13288 23000 13290
rect 21265 13232 21270 13288
rect 21326 13232 23000 13288
rect 21265 13230 23000 13232
rect 19977 13227 20043 13230
rect 21265 13227 21331 13230
rect 22200 13200 23000 13230
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 21265 12882 21331 12885
rect 22200 12882 23000 12912
rect 21265 12880 23000 12882
rect 21265 12824 21270 12880
rect 21326 12824 23000 12880
rect 21265 12822 23000 12824
rect 21265 12819 21331 12822
rect 22200 12792 23000 12822
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 22200 12474 23000 12504
rect 19566 12414 23000 12474
rect 19149 12338 19215 12341
rect 19566 12338 19626 12414
rect 22200 12384 23000 12414
rect 19149 12336 19626 12338
rect 19149 12280 19154 12336
rect 19210 12280 19626 12336
rect 19149 12278 19626 12280
rect 19149 12275 19215 12278
rect 20253 12202 20319 12205
rect 20253 12200 22202 12202
rect 20253 12144 20258 12200
rect 20314 12144 22202 12200
rect 20253 12142 22202 12144
rect 20253 12139 20319 12142
rect 22142 12096 22202 12142
rect 22142 12006 23000 12096
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 16941 11794 17007 11797
rect 17350 11794 17356 11796
rect 16941 11792 17356 11794
rect 16941 11736 16946 11792
rect 17002 11736 17356 11792
rect 16941 11734 17356 11736
rect 16941 11731 17007 11734
rect 17350 11732 17356 11734
rect 17420 11732 17426 11796
rect 21725 11658 21791 11661
rect 22200 11658 23000 11688
rect 21725 11656 23000 11658
rect 21725 11600 21730 11656
rect 21786 11600 23000 11656
rect 21725 11598 23000 11600
rect 21725 11595 21791 11598
rect 22200 11568 23000 11598
rect 0 11522 800 11552
rect 1485 11522 1551 11525
rect 0 11520 1551 11522
rect 0 11464 1490 11520
rect 1546 11464 1551 11520
rect 0 11462 1551 11464
rect 0 11432 800 11462
rect 1485 11459 1551 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 13537 11250 13603 11253
rect 19977 11250 20043 11253
rect 13537 11248 20043 11250
rect 13537 11192 13542 11248
rect 13598 11192 19982 11248
rect 20038 11192 20043 11248
rect 13537 11190 20043 11192
rect 13537 11187 13603 11190
rect 19977 11187 20043 11190
rect 21449 11250 21515 11253
rect 22200 11250 23000 11280
rect 21449 11248 23000 11250
rect 21449 11192 21454 11248
rect 21510 11192 23000 11248
rect 21449 11190 23000 11192
rect 21449 11187 21515 11190
rect 22200 11160 23000 11190
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 22200 10842 23000 10872
rect 22142 10752 23000 10842
rect 17953 10706 18019 10709
rect 22142 10706 22202 10752
rect 17953 10704 22202 10706
rect 17953 10648 17958 10704
rect 18014 10648 22202 10704
rect 17953 10646 22202 10648
rect 17953 10643 18019 10646
rect 21357 10434 21423 10437
rect 22200 10434 23000 10464
rect 21357 10432 23000 10434
rect 21357 10376 21362 10432
rect 21418 10376 23000 10432
rect 21357 10374 23000 10376
rect 21357 10371 21423 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 22200 10344 23000 10374
rect 19139 10303 19455 10304
rect 18229 10026 18295 10029
rect 22200 10026 23000 10056
rect 18229 10024 23000 10026
rect 18229 9968 18234 10024
rect 18290 9968 23000 10024
rect 18229 9966 23000 9968
rect 18229 9963 18295 9966
rect 22200 9936 23000 9966
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 17769 9754 17835 9757
rect 17726 9752 17835 9754
rect 17726 9696 17774 9752
rect 17830 9696 17835 9752
rect 17726 9691 17835 9696
rect 17726 9346 17786 9691
rect 21449 9618 21515 9621
rect 22200 9618 23000 9648
rect 21449 9616 23000 9618
rect 21449 9560 21454 9616
rect 21510 9560 23000 9616
rect 21449 9558 23000 9560
rect 21449 9555 21515 9558
rect 22200 9528 23000 9558
rect 17861 9346 17927 9349
rect 17726 9344 17927 9346
rect 17726 9288 17866 9344
rect 17922 9288 17927 9344
rect 17726 9286 17927 9288
rect 17861 9283 17927 9286
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 22200 9210 23000 9240
rect 19566 9150 23000 9210
rect 19241 9074 19307 9077
rect 19566 9074 19626 9150
rect 22200 9120 23000 9150
rect 19241 9072 19626 9074
rect 19241 9016 19246 9072
rect 19302 9016 19626 9072
rect 19241 9014 19626 9016
rect 19241 9011 19307 9014
rect 18965 8938 19031 8941
rect 18965 8936 22202 8938
rect 18965 8880 18970 8936
rect 19026 8880 22202 8936
rect 18965 8878 22202 8880
rect 18965 8875 19031 8878
rect 22142 8832 22202 8878
rect 22142 8742 23000 8832
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 18505 8666 18571 8669
rect 19006 8666 19012 8668
rect 18505 8664 19012 8666
rect 18505 8608 18510 8664
rect 18566 8608 19012 8664
rect 18505 8606 19012 8608
rect 18505 8603 18571 8606
rect 19006 8604 19012 8606
rect 19076 8604 19082 8668
rect 14549 8394 14615 8397
rect 18689 8394 18755 8397
rect 14549 8392 18755 8394
rect 14549 8336 14554 8392
rect 14610 8336 18694 8392
rect 18750 8336 18755 8392
rect 14549 8334 18755 8336
rect 14549 8331 14615 8334
rect 18689 8331 18755 8334
rect 18965 8394 19031 8397
rect 22200 8394 23000 8424
rect 18965 8392 23000 8394
rect 18965 8336 18970 8392
rect 19026 8336 23000 8392
rect 18965 8334 23000 8336
rect 18965 8331 19031 8334
rect 22200 8304 23000 8334
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 17953 7986 18019 7989
rect 22200 7986 23000 8016
rect 17953 7984 23000 7986
rect 17953 7928 17958 7984
rect 18014 7928 23000 7984
rect 17953 7926 23000 7928
rect 17953 7923 18019 7926
rect 22200 7896 23000 7926
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 22200 7578 23000 7608
rect 22142 7488 23000 7578
rect 17861 7442 17927 7445
rect 19701 7442 19767 7445
rect 17861 7440 19767 7442
rect 17861 7384 17866 7440
rect 17922 7384 19706 7440
rect 19762 7384 19767 7440
rect 17861 7382 19767 7384
rect 17861 7379 17927 7382
rect 19701 7379 19767 7382
rect 20345 7442 20411 7445
rect 22142 7442 22202 7488
rect 20345 7440 22202 7442
rect 20345 7384 20350 7440
rect 20406 7384 22202 7440
rect 20345 7382 22202 7384
rect 20345 7379 20411 7382
rect 18321 7306 18387 7309
rect 18321 7304 19626 7306
rect 18321 7248 18326 7304
rect 18382 7248 19626 7304
rect 18321 7246 19626 7248
rect 18321 7243 18387 7246
rect 19566 7170 19626 7246
rect 22200 7170 23000 7200
rect 19566 7110 23000 7170
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 22200 7080 23000 7110
rect 19139 7039 19455 7040
rect 18965 6762 19031 6765
rect 21357 6762 21423 6765
rect 22200 6762 23000 6792
rect 18965 6760 23000 6762
rect 18965 6704 18970 6760
rect 19026 6704 21362 6760
rect 21418 6704 23000 6760
rect 18965 6702 23000 6704
rect 18965 6699 19031 6702
rect 21357 6699 21423 6702
rect 22200 6672 23000 6702
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 20805 6490 20871 6493
rect 18094 6488 20871 6490
rect 18094 6432 20810 6488
rect 20866 6432 20871 6488
rect 18094 6430 20871 6432
rect 9765 6354 9831 6357
rect 18094 6354 18154 6430
rect 20805 6427 20871 6430
rect 9765 6352 18154 6354
rect 9765 6296 9770 6352
rect 9826 6296 18154 6352
rect 9765 6294 18154 6296
rect 18321 6354 18387 6357
rect 22200 6354 23000 6384
rect 18321 6352 23000 6354
rect 18321 6296 18326 6352
rect 18382 6296 23000 6352
rect 18321 6294 23000 6296
rect 9765 6291 9831 6294
rect 18321 6291 18387 6294
rect 22200 6264 23000 6294
rect 17953 6218 18019 6221
rect 17953 6216 19626 6218
rect 17953 6160 17958 6216
rect 18014 6160 19626 6216
rect 17953 6158 19626 6160
rect 17953 6155 18019 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 19566 5946 19626 6158
rect 22200 5946 23000 5976
rect 19566 5886 23000 5946
rect 22200 5856 23000 5886
rect 18454 5612 18460 5676
rect 18524 5674 18530 5676
rect 19517 5674 19583 5677
rect 18524 5672 19583 5674
rect 18524 5616 19522 5672
rect 19578 5616 19583 5672
rect 18524 5614 19583 5616
rect 18524 5612 18530 5614
rect 19517 5611 19583 5614
rect 21590 5614 22202 5674
rect 17953 5538 18019 5541
rect 21590 5538 21650 5614
rect 17953 5536 21650 5538
rect 17953 5480 17958 5536
rect 18014 5480 21650 5536
rect 17953 5478 21650 5480
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 17953 5475 18019 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 17309 5404 17375 5405
rect 17309 5402 17356 5404
rect 17264 5400 17356 5402
rect 17264 5344 17314 5400
rect 17264 5342 17356 5344
rect 17309 5340 17356 5342
rect 17420 5340 17426 5404
rect 17309 5339 17375 5340
rect 18045 5130 18111 5133
rect 22200 5130 23000 5160
rect 18045 5128 23000 5130
rect 18045 5072 18050 5128
rect 18106 5072 23000 5128
rect 18045 5070 23000 5072
rect 18045 5067 18111 5070
rect 22200 5040 23000 5070
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 17861 4722 17927 4725
rect 22200 4722 23000 4752
rect 17861 4720 23000 4722
rect 17861 4664 17866 4720
rect 17922 4664 23000 4720
rect 17861 4662 23000 4664
rect 17861 4659 17927 4662
rect 22200 4632 23000 4662
rect 8569 4586 8635 4589
rect 19609 4586 19675 4589
rect 8569 4584 19675 4586
rect 8569 4528 8574 4584
rect 8630 4528 19614 4584
rect 19670 4528 19675 4584
rect 8569 4526 19675 4528
rect 8569 4523 8635 4526
rect 19609 4523 19675 4526
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 22200 4314 23000 4344
rect 22142 4224 23000 4314
rect 16481 4178 16547 4181
rect 17309 4178 17375 4181
rect 16481 4176 17375 4178
rect 16481 4120 16486 4176
rect 16542 4120 17314 4176
rect 17370 4120 17375 4176
rect 16481 4118 17375 4120
rect 16481 4115 16547 4118
rect 17309 4115 17375 4118
rect 17953 4178 18019 4181
rect 22142 4178 22202 4224
rect 17953 4176 22202 4178
rect 17953 4120 17958 4176
rect 18014 4120 22202 4176
rect 17953 4118 22202 4120
rect 17953 4115 18019 4118
rect 13353 4042 13419 4045
rect 19977 4042 20043 4045
rect 13353 4040 20043 4042
rect 13353 3984 13358 4040
rect 13414 3984 19982 4040
rect 20038 3984 20043 4040
rect 13353 3982 20043 3984
rect 13353 3979 13419 3982
rect 19977 3979 20043 3982
rect 20529 3906 20595 3909
rect 22200 3906 23000 3936
rect 20529 3904 23000 3906
rect 20529 3848 20534 3904
rect 20590 3848 23000 3904
rect 20529 3846 23000 3848
rect 20529 3843 20595 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 18229 3636 18295 3637
rect 18229 3634 18276 3636
rect 18184 3632 18276 3634
rect 18184 3576 18234 3632
rect 18184 3574 18276 3576
rect 18229 3572 18276 3574
rect 18340 3572 18346 3636
rect 18229 3571 18295 3572
rect 13261 3498 13327 3501
rect 18597 3498 18663 3501
rect 13261 3496 18663 3498
rect 13261 3440 13266 3496
rect 13322 3440 18602 3496
rect 18658 3440 18663 3496
rect 13261 3438 18663 3440
rect 13261 3435 13327 3438
rect 18597 3435 18663 3438
rect 18781 3498 18847 3501
rect 22200 3498 23000 3528
rect 18781 3496 23000 3498
rect 18781 3440 18786 3496
rect 18842 3440 23000 3496
rect 18781 3438 23000 3440
rect 18781 3435 18847 3438
rect 22200 3408 23000 3438
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 14549 3090 14615 3093
rect 19333 3090 19399 3093
rect 14549 3088 19399 3090
rect 14549 3032 14554 3088
rect 14610 3032 19338 3088
rect 19394 3032 19399 3088
rect 14549 3030 19399 3032
rect 14549 3027 14615 3030
rect 19333 3027 19399 3030
rect 20529 3090 20595 3093
rect 22200 3090 23000 3120
rect 20529 3088 23000 3090
rect 20529 3032 20534 3088
rect 20590 3032 23000 3088
rect 20529 3030 23000 3032
rect 20529 3027 20595 3030
rect 22200 3000 23000 3030
rect 14825 2954 14891 2957
rect 19885 2954 19951 2957
rect 14825 2952 19951 2954
rect 14825 2896 14830 2952
rect 14886 2896 19890 2952
rect 19946 2896 19951 2952
rect 14825 2894 19951 2896
rect 14825 2891 14891 2894
rect 19885 2891 19951 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 20529 2682 20595 2685
rect 22200 2682 23000 2712
rect 20529 2680 23000 2682
rect 20529 2624 20534 2680
rect 20590 2624 23000 2680
rect 20529 2622 23000 2624
rect 20529 2619 20595 2622
rect 22200 2592 23000 2622
rect 20529 2410 20595 2413
rect 20529 2408 22202 2410
rect 20529 2352 20534 2408
rect 20590 2352 22202 2408
rect 20529 2350 22202 2352
rect 20529 2347 20595 2350
rect 22142 2304 22202 2350
rect 22142 2214 23000 2304
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 20253 1866 20319 1869
rect 22200 1866 23000 1896
rect 20253 1864 23000 1866
rect 20253 1808 20258 1864
rect 20314 1808 23000 1864
rect 20253 1806 23000 1808
rect 20253 1803 20319 1806
rect 22200 1776 23000 1806
rect 19241 1458 19307 1461
rect 22200 1458 23000 1488
rect 19241 1456 23000 1458
rect 19241 1400 19246 1456
rect 19302 1400 23000 1456
rect 19241 1398 23000 1400
rect 19241 1395 19307 1398
rect 22200 1368 23000 1398
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 18276 15948 18340 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 17356 14316 17420 14380
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 18460 13968 18524 13972
rect 18460 13912 18474 13968
rect 18474 13912 18524 13968
rect 18460 13908 18524 13912
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 19012 13424 19076 13428
rect 19012 13368 19026 13424
rect 19026 13368 19076 13424
rect 19012 13364 19076 13368
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 17356 11732 17420 11796
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 19012 8604 19076 8668
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 18460 5612 18524 5676
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 17356 5400 17420 5404
rect 17356 5344 17370 5400
rect 17370 5344 17420 5400
rect 17356 5340 17420 5344
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 18276 3632 18340 3636
rect 18276 3576 18290 3632
rect 18290 3576 18340 3632
rect 18276 3572 18340 3576
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 18275 16012 18341 16013
rect 18275 15948 18276 16012
rect 18340 15948 18341 16012
rect 18275 15947 18341 15948
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 17355 14380 17421 14381
rect 17355 14316 17356 14380
rect 17420 14316 17421 14380
rect 17355 14315 17421 14316
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 17358 11797 17418 14315
rect 17355 11796 17421 11797
rect 17355 11732 17356 11796
rect 17420 11732 17421 11796
rect 17355 11731 17421 11732
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 17358 5405 17418 11731
rect 17355 5404 17421 5405
rect 17355 5340 17356 5404
rect 17420 5340 17421 5404
rect 17355 5339 17421 5340
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 18278 3637 18338 15947
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 18459 13972 18525 13973
rect 18459 13908 18460 13972
rect 18524 13908 18525 13972
rect 18459 13907 18525 13908
rect 18462 5677 18522 13907
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19011 13428 19077 13429
rect 19011 13364 19012 13428
rect 19076 13364 19077 13428
rect 19011 13363 19077 13364
rect 19014 8669 19074 13363
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19011 8668 19077 8669
rect 19011 8604 19012 8668
rect 19076 8604 19077 8668
rect 19011 8603 19077 8604
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 18459 5676 18525 5677
rect 18459 5612 18460 5676
rect 18524 5612 18525 5676
rect 18459 5611 18525 5612
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 18275 3636 18341 3637
rect 18275 3572 18276 3636
rect 18340 3572 18341 3636
rect 18275 3571 18341 3572
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 19780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 17020 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 16100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 17940 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 17296 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 2392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 7360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 10948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 4876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 5796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 13340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15364 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17940 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12972 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 20424 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 15180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 14812 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1649977179
transform 1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_130
timestamp 1649977179
transform 1 0 13064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_14
timestamp 1649977179
transform 1 0 2392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_38
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_41
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_46
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_64
timestamp 1649977179
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1649977179
transform 1 0 7360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1649977179
transform 1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_97
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1649977179
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_115
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1649977179
transform 1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_160
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1649977179
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp 1649977179
transform 1 0 17572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1649977179
transform 1 0 18584 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_202
timestamp 1649977179
transform 1 0 19688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1649977179
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1649977179
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1649977179
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_36
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_48
timestamp 1649977179
transform 1 0 5520 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_60
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_72
timestamp 1649977179
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 1649977179
transform 1 0 14628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_152
timestamp 1649977179
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_161
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1649977179
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_156
timestamp 1649977179
transform 1 0 15456 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_191
timestamp 1649977179
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1649977179
transform 1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1649977179
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_159
timestamp 1649977179
transform 1 0 15732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_170
timestamp 1649977179
transform 1 0 16744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1649977179
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_184
timestamp 1649977179
transform 1 0 18032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1649977179
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_183
timestamp 1649977179
transform 1 0 17940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1649977179
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1649977179
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1649977179
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1649977179
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_173
timestamp 1649977179
transform 1 0 17020 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_183
timestamp 1649977179
transform 1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_194
timestamp 1649977179
transform 1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_198
timestamp 1649977179
transform 1 0 19320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_202
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_207
timestamp 1649977179
transform 1 0 20148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_218
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_222
timestamp 1649977179
transform 1 0 21528 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_169
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_217
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1649977179
transform 1 0 17204 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1649977179
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_183
timestamp 1649977179
transform 1 0 17940 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1649977179
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_199
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_203
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1649977179
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_174
timestamp 1649977179
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1649977179
transform 1 0 20148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1649977179
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1649977179
transform 1 0 21528 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1649977179
transform 1 0 17296 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1649977179
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_196
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1649977179
transform 1 0 19504 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_211
timestamp 1649977179
transform 1 0 20516 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1649977179
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_162
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1649977179
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_199
timestamp 1649977179
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_204
timestamp 1649977179
transform 1 0 19872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_141
timestamp 1649977179
transform 1 0 14076 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1649977179
transform 1 0 18032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_195
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_199
timestamp 1649977179
transform 1 0 19412 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_164
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1649977179
transform 1 0 17756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1649977179
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1649977179
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1649977179
transform 1 0 21528 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_186
timestamp 1649977179
transform 1 0 18216 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1649977179
transform 1 0 18676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_202
timestamp 1649977179
transform 1 0 19688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1649977179
transform 1 0 20608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1649977179
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_211
timestamp 1649977179
transform 1 0 20516 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_216
timestamp 1649977179
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1649977179
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1649977179
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_160
timestamp 1649977179
transform 1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_172
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_195
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1649977179
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_211
timestamp 1649977179
transform 1 0 20516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_108
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_116
timestamp 1649977179
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1649977179
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1649977179
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1649977179
transform 1 0 20424 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1649977179
transform 1 0 20884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_141
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1649977179
transform 1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_171
timestamp 1649977179
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_182
timestamp 1649977179
transform 1 0 17848 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1649977179
transform 1 0 20424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1649977179
transform 1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_171
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_203
timestamp 1649977179
transform 1 0 19780 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_87
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1649977179
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1649977179
transform 1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_138
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_150
timestamp 1649977179
transform 1 0 14904 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_187
timestamp 1649977179
transform 1 0 18308 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1649977179
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_179
timestamp 1649977179
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1649977179
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_145
timestamp 1649977179
transform 1 0 14444 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1649977179
transform 1 0 16008 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1649977179
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_105
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_124
timestamp 1649977179
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1649977179
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_175
timestamp 1649977179
transform 1 0 17204 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_179
timestamp 1649977179
transform 1 0 17572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_183
timestamp 1649977179
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_191
timestamp 1649977179
transform 1 0 18676 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_138
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_150
timestamp 1649977179
transform 1 0 14904 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_158
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_196
timestamp 1649977179
transform 1 0 19136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_202
timestamp 1649977179
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1649977179
transform 1 0 17756 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_185
timestamp 1649977179
transform 1 0 18124 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_117
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1649977179
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_139
timestamp 1649977179
transform 1 0 13892 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1649977179
transform 1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1649977179
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_161
timestamp 1649977179
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1649977179
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_135
timestamp 1649977179
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_139
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_145
timestamp 1649977179
transform 1 0 14444 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1649977179
transform 1 0 14720 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_191
timestamp 1649977179
transform 1 0 18676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1649977179
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_92
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_111
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_129
timestamp 1649977179
transform 1 0 12972 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_159
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_181
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1649977179
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_88
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_115
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_141
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1649977179
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1649977179
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_94
timestamp 1649977179
transform 1 0 9752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1649977179
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_110
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1649977179
transform 1 0 13156 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_147
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_160
timestamp 1649977179
transform 1 0 15824 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_168
timestamp 1649977179
transform 1 0 16560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1649977179
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_71
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_89
timestamp 1649977179
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_94
timestamp 1649977179
transform 1 0 9752 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1649977179
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1649977179
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_133
timestamp 1649977179
transform 1 0 13340 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_176
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_182
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1649977179
transform 1 0 18400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _48_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform 1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 19688 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 16560 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 14996 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 13616 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform 1 0 18952 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform -1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform -1 0 16376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform -1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform 1 0 18768 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1649977179
transform -1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1649977179
transform -1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1649977179
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp 1649977179
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _88_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 16376 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 19780 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 20240 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 17664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 18952 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 18952 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1649977179
transform 1 0 20516 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform -1 0 20148 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18860 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14260 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17388 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18676 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15916 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18492 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17940 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11960 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12512 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14260 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15916 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16836 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13248 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11960 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_0__108 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_0__110
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18216 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_0__109
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20148 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 20240 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 20332 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_1__112
timestamp 1649977179
transform -1 0 18952 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19872 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_1__118
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18676 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 19412 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 20792 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20424 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20884 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_1__105
timestamp 1649977179
transform -1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_6.mux_l2_in_1__106
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l1_in_1__107
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18032 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18768 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_10.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14996 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_12.mux_l2_in_0__114
timestamp 1649977179
transform 1 0 15272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15640 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_14.mux_l2_in_0__115
timestamp 1649977179
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15640 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_0__116
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15364 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_18.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19780 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8740 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_20.mux_l2_in_0__95
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20516 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_22.mux_l2_in_0__96
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_1__97
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17756 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_26.mux_l2_in_0__98
timestamp 1649977179
transform 1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17112 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_28.mux_l2_in_0__99
timestamp 1649977179
transform -1 0 7636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_30.mux_l2_in_0__100
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_0__101
timestamp 1649977179
transform 1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8648 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_34.mux_l2_in_0__102
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_36.mux_l2_in_0__103
timestamp 1649977179
transform -1 0 8188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18676 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_38.mux_l2_in_0__104
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 19412 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 18032 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 20516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 19780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
<< labels >>
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 SC_IN_TOP
port 0 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_1_
port 4 nsew signal input
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 ccff_head
port 5 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 ccff_tail
port 6 nsew signal tristate
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 7 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 8 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 9 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 10 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 11 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 12 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 13 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 14 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 15 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 16 nsew signal input
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 17 nsew signal input
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 18 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 19 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 20 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 21 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 22 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 23 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 24 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 25 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 26 nsew signal input
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 27 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 28 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 29 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 30 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 31 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 32 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 33 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 34 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 35 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 36 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 37 nsew signal tristate
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 38 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 39 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 40 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 41 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 42 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 43 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 44 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 45 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 46 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 47 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 48 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 49 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 50 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 51 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 52 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 53 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 54 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 55 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 56 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 57 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 58 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 59 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 60 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 61 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 62 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 63 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 64 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 65 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 66 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 67 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 68 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 69 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 70 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 71 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 72 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 73 nsew signal tristate
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 74 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 75 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 76 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 77 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 78 nsew signal tristate
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 79 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 80 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 81 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 82 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 83 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 84 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 85 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 86 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 87 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 88 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 89 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 90 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 91 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 92 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 93 nsew signal input
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 94 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 95 nsew signal input
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 right_top_grid_pin_1_
port 96 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
