magic
tech sky130A
magscale 1 2
timestamp 1679357491
<< viali >>
rect 15485 24361 15519 24395
rect 17601 24361 17635 24395
rect 18153 24293 18187 24327
rect 23765 24293 23799 24327
rect 3249 24225 3283 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 12817 24225 12851 24259
rect 16221 24225 16255 24259
rect 16405 24225 16439 24259
rect 18797 24225 18831 24259
rect 20085 24225 20119 24259
rect 20821 24225 20855 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9321 24157 9355 24191
rect 9781 24157 9815 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 16957 24157 16991 24191
rect 18521 24157 18555 24191
rect 19809 24157 19843 24191
rect 21097 24157 21131 24191
rect 22017 24157 22051 24191
rect 24961 24157 24995 24191
rect 5825 24089 5859 24123
rect 14381 24089 14415 24123
rect 15393 24089 15427 24123
rect 16773 24089 16807 24123
rect 22845 24089 22879 24123
rect 3985 24021 4019 24055
rect 6561 24021 6595 24055
rect 9137 24021 9171 24055
rect 14473 24021 14507 24055
rect 15761 24021 15795 24055
rect 16129 24021 16163 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 19901 24021 19935 24055
rect 20637 24021 20671 24055
rect 24593 24021 24627 24055
rect 25053 24021 25087 24055
rect 16865 23817 16899 23851
rect 3985 23749 4019 23783
rect 5825 23749 5859 23783
rect 9137 23749 9171 23783
rect 10885 23749 10919 23783
rect 14473 23749 14507 23783
rect 17233 23749 17267 23783
rect 25145 23749 25179 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6561 23681 6595 23715
rect 7941 23681 7975 23715
rect 9781 23681 9815 23715
rect 12081 23681 12115 23715
rect 14381 23681 14415 23715
rect 15945 23681 15979 23715
rect 20177 23681 20211 23715
rect 20637 23681 20671 23715
rect 22017 23681 22051 23715
rect 6837 23613 6871 23647
rect 12541 23613 12575 23647
rect 14565 23613 14599 23647
rect 16037 23613 16071 23647
rect 16221 23613 16255 23647
rect 17325 23613 17359 23647
rect 17509 23613 17543 23647
rect 17877 23613 17911 23647
rect 18153 23613 18187 23647
rect 20913 23613 20947 23647
rect 22109 23613 22143 23647
rect 22385 23613 22419 23647
rect 23857 23613 23891 23647
rect 14013 23545 14047 23579
rect 15577 23545 15611 23579
rect 1777 23477 1811 23511
rect 19625 23477 19659 23511
rect 21833 23477 21867 23511
rect 25237 23477 25271 23511
rect 18889 23273 18923 23307
rect 21189 23273 21223 23307
rect 3249 23137 3283 23171
rect 6561 23137 6595 23171
rect 8217 23137 8251 23171
rect 10517 23137 10551 23171
rect 12173 23137 12207 23171
rect 14933 23137 14967 23171
rect 15209 23137 15243 23171
rect 17141 23137 17175 23171
rect 19441 23137 19475 23171
rect 21557 23137 21591 23171
rect 21833 23137 21867 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 3985 23069 4019 23103
rect 4261 23069 4295 23103
rect 5549 23069 5583 23103
rect 7205 23069 7239 23103
rect 9413 23069 9447 23103
rect 9873 23069 9907 23103
rect 11713 23069 11747 23103
rect 13737 23069 13771 23103
rect 14473 23069 14507 23103
rect 21465 23069 21499 23103
rect 24961 23069 24995 23103
rect 17424 23001 17458 23035
rect 19717 23001 19751 23035
rect 23765 23001 23799 23035
rect 9229 22933 9263 22967
rect 13553 22933 13587 22967
rect 16681 22933 16715 22967
rect 23305 22933 23339 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 11713 22729 11747 22763
rect 12173 22729 12207 22763
rect 15301 22729 15335 22763
rect 15945 22729 15979 22763
rect 17049 22729 17083 22763
rect 17233 22729 17267 22763
rect 18981 22729 19015 22763
rect 20177 22729 20211 22763
rect 22385 22729 22419 22763
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 8769 22661 8803 22695
rect 13829 22661 13863 22695
rect 17601 22661 17635 22695
rect 1685 22593 1719 22627
rect 2973 22593 3007 22627
rect 4813 22593 4847 22627
rect 6653 22593 6687 22627
rect 7573 22593 7607 22627
rect 12081 22593 12115 22627
rect 13093 22593 13127 22627
rect 13553 22593 13587 22627
rect 15853 22593 15887 22627
rect 16957 22593 16991 22627
rect 18521 22593 18555 22627
rect 19349 22593 19383 22627
rect 20545 22593 20579 22627
rect 24501 22593 24535 22627
rect 9413 22525 9447 22559
rect 9689 22525 9723 22559
rect 12265 22525 12299 22559
rect 17693 22525 17727 22559
rect 17785 22525 17819 22559
rect 19441 22525 19475 22559
rect 19625 22525 19659 22559
rect 20637 22525 20671 22559
rect 20729 22525 20763 22559
rect 22477 22525 22511 22559
rect 22661 22525 22695 22559
rect 24593 22525 24627 22559
rect 24685 22525 24719 22559
rect 1869 22457 1903 22491
rect 11161 22457 11195 22491
rect 21649 22457 21683 22491
rect 6745 22389 6779 22423
rect 12909 22389 12943 22423
rect 22017 22389 22051 22423
rect 23673 22389 23707 22423
rect 24133 22389 24167 22423
rect 9965 22185 9999 22219
rect 10872 22185 10906 22219
rect 14841 22117 14875 22151
rect 17325 22117 17359 22151
rect 2881 22049 2915 22083
rect 6101 22049 6135 22083
rect 8309 22049 8343 22083
rect 12357 22049 12391 22083
rect 16589 22049 16623 22083
rect 17969 22049 18003 22083
rect 20085 22049 20119 22083
rect 20453 22049 20487 22083
rect 22201 22049 22235 22083
rect 22477 22049 22511 22083
rect 25237 22049 25271 22083
rect 2237 21981 2271 22015
rect 4077 21981 4111 22015
rect 4905 21981 4939 22015
rect 5549 21981 5583 22015
rect 7389 21981 7423 22015
rect 9505 21981 9539 22015
rect 10149 21981 10183 22015
rect 10609 21981 10643 22015
rect 13553 21981 13587 22015
rect 17785 21981 17819 22015
rect 19809 21981 19843 22015
rect 22753 21981 22787 22015
rect 4261 21913 4295 21947
rect 14657 21913 14691 21947
rect 15393 21913 15427 21947
rect 18613 21913 18647 21947
rect 20729 21913 20763 21947
rect 25053 21913 25087 21947
rect 4721 21845 4755 21879
rect 9321 21845 9355 21879
rect 15485 21845 15519 21879
rect 16037 21845 16071 21879
rect 16405 21845 16439 21879
rect 16497 21845 16531 21879
rect 17693 21845 17727 21879
rect 18705 21845 18739 21879
rect 19441 21845 19475 21879
rect 19901 21845 19935 21879
rect 23765 21845 23799 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 12081 21641 12115 21675
rect 12449 21641 12483 21675
rect 15485 21641 15519 21675
rect 19993 21641 20027 21675
rect 24041 21641 24075 21675
rect 25053 21641 25087 21675
rect 1685 21573 1719 21607
rect 13553 21573 13587 21607
rect 17509 21573 17543 21607
rect 2973 21505 3007 21539
rect 4813 21505 4847 21539
rect 7481 21505 7515 21539
rect 15853 21505 15887 21539
rect 17417 21505 17451 21539
rect 18245 21505 18279 21539
rect 20821 21505 20855 21539
rect 24961 21505 24995 21539
rect 1869 21437 1903 21471
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 7757 21437 7791 21471
rect 9137 21437 9171 21471
rect 9413 21437 9447 21471
rect 12541 21437 12575 21471
rect 12633 21437 12667 21471
rect 13277 21437 13311 21471
rect 15945 21437 15979 21471
rect 16129 21437 16163 21471
rect 17693 21437 17727 21471
rect 18521 21437 18555 21471
rect 20913 21437 20947 21471
rect 21097 21437 21131 21471
rect 22293 21437 22327 21471
rect 24317 21437 24351 21471
rect 25145 21437 25179 21471
rect 6837 21301 6871 21335
rect 10885 21301 10919 21335
rect 15025 21301 15059 21335
rect 17049 21301 17083 21335
rect 20453 21301 20487 21335
rect 22556 21301 22590 21335
rect 24593 21301 24627 21335
rect 12909 21097 12943 21131
rect 15485 21097 15519 21131
rect 16865 21097 16899 21131
rect 19625 21097 19659 21131
rect 24225 21097 24259 21131
rect 14289 21029 14323 21063
rect 17509 21029 17543 21063
rect 22109 21029 22143 21063
rect 2881 20961 2915 20995
rect 4445 20961 4479 20995
rect 7389 20961 7423 20995
rect 10425 20961 10459 20995
rect 10609 20961 10643 20995
rect 11161 20961 11195 20995
rect 14749 20961 14783 20995
rect 14933 20961 14967 20995
rect 16037 20961 16071 20995
rect 18061 20961 18095 20995
rect 20361 20961 20395 20995
rect 20637 20961 20671 20995
rect 22753 20961 22787 20995
rect 24961 20961 24995 20995
rect 2237 20893 2271 20927
rect 4077 20893 4111 20927
rect 6009 20893 6043 20927
rect 7113 20893 7147 20927
rect 9321 20893 9355 20927
rect 13553 20893 13587 20927
rect 14657 20893 14691 20927
rect 18889 20893 18923 20927
rect 22477 20893 22511 20927
rect 24777 20893 24811 20927
rect 11437 20825 11471 20859
rect 16773 20825 16807 20859
rect 17969 20825 18003 20859
rect 24869 20825 24903 20859
rect 5825 20757 5859 20791
rect 9137 20757 9171 20791
rect 9965 20757 9999 20791
rect 10333 20757 10367 20791
rect 15853 20757 15887 20791
rect 15945 20757 15979 20791
rect 17877 20757 17911 20791
rect 24409 20757 24443 20791
rect 12449 20553 12483 20587
rect 15945 20553 15979 20587
rect 18705 20553 18739 20587
rect 22385 20553 22419 20587
rect 22477 20553 22511 20587
rect 23213 20485 23247 20519
rect 1869 20417 1903 20451
rect 2973 20417 3007 20451
rect 6009 20417 6043 20451
rect 7113 20417 7147 20451
rect 8585 20417 8619 20451
rect 13553 20417 13587 20451
rect 15853 20417 15887 20451
rect 19257 20417 19291 20451
rect 1593 20349 1627 20383
rect 3341 20349 3375 20383
rect 7389 20349 7423 20383
rect 9045 20349 9079 20383
rect 9321 20349 9355 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 13829 20349 13863 20383
rect 16957 20349 16991 20383
rect 17233 20349 17267 20383
rect 19533 20349 19567 20383
rect 21005 20349 21039 20383
rect 22569 20349 22603 20383
rect 23489 20349 23523 20383
rect 23765 20349 23799 20383
rect 4721 20281 4755 20315
rect 5365 20281 5399 20315
rect 12081 20281 12115 20315
rect 5825 20213 5859 20247
rect 8401 20213 8435 20247
rect 10793 20213 10827 20247
rect 15301 20213 15335 20247
rect 22017 20213 22051 20247
rect 25237 20213 25271 20247
rect 6469 20009 6503 20043
rect 14933 20009 14967 20043
rect 17693 20009 17727 20043
rect 7113 19941 7147 19975
rect 13369 19941 13403 19975
rect 16313 19941 16347 19975
rect 22845 19941 22879 19975
rect 2881 19873 2915 19907
rect 4813 19873 4847 19907
rect 9781 19873 9815 19907
rect 10977 19873 11011 19907
rect 11621 19873 11655 19907
rect 15485 19873 15519 19907
rect 16865 19873 16899 19907
rect 18245 19873 18279 19907
rect 19993 19873 20027 19907
rect 21097 19873 21131 19907
rect 25145 19873 25179 19907
rect 2237 19805 2271 19839
rect 4537 19805 4571 19839
rect 6009 19805 6043 19839
rect 6653 19805 6687 19839
rect 7297 19805 7331 19839
rect 7941 19805 7975 19839
rect 8585 19805 8619 19839
rect 9597 19805 9631 19839
rect 9689 19805 9723 19839
rect 14473 19805 14507 19839
rect 19809 19805 19843 19839
rect 24961 19805 24995 19839
rect 11897 19737 11931 19771
rect 15301 19737 15335 19771
rect 15393 19737 15427 19771
rect 16681 19737 16715 19771
rect 18153 19737 18187 19771
rect 21373 19737 21407 19771
rect 25053 19737 25087 19771
rect 5825 19669 5859 19703
rect 7757 19669 7791 19703
rect 9229 19669 9263 19703
rect 10425 19669 10459 19703
rect 10793 19669 10827 19703
rect 10885 19669 10919 19703
rect 14289 19669 14323 19703
rect 16773 19669 16807 19703
rect 18061 19669 18095 19703
rect 19441 19669 19475 19703
rect 19901 19669 19935 19703
rect 23765 19669 23799 19703
rect 24593 19669 24627 19703
rect 4169 19465 4203 19499
rect 5457 19465 5491 19499
rect 6561 19465 6595 19499
rect 7757 19465 7791 19499
rect 10885 19465 10919 19499
rect 14473 19465 14507 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 20361 19465 20395 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 22477 19465 22511 19499
rect 25145 19465 25179 19499
rect 19533 19397 19567 19431
rect 1961 19329 1995 19363
rect 4353 19329 4387 19363
rect 5641 19329 5675 19363
rect 6009 19329 6043 19363
rect 6745 19329 6779 19363
rect 7389 19329 7423 19363
rect 7941 19329 7975 19363
rect 8217 19329 8251 19363
rect 12081 19329 12115 19363
rect 12725 19329 12759 19363
rect 16313 19329 16347 19363
rect 16957 19329 16991 19363
rect 19625 19329 19659 19363
rect 20729 19329 20763 19363
rect 2237 19261 2271 19295
rect 9137 19261 9171 19295
rect 9413 19261 9447 19295
rect 13001 19261 13035 19295
rect 15393 19261 15427 19295
rect 15577 19261 15611 19295
rect 17233 19261 17267 19295
rect 18705 19261 18739 19295
rect 19717 19261 19751 19295
rect 20821 19261 20855 19295
rect 21005 19261 21039 19295
rect 22569 19261 22603 19295
rect 23397 19261 23431 19295
rect 23673 19261 23707 19295
rect 5365 19193 5399 19227
rect 7205 19193 7239 19227
rect 4077 19125 4111 19159
rect 4721 19125 4755 19159
rect 5825 19125 5859 19159
rect 8033 19125 8067 19159
rect 8677 19125 8711 19159
rect 12173 19125 12207 19159
rect 16129 19125 16163 19159
rect 19165 19125 19199 19159
rect 23213 19125 23247 19159
rect 1961 18921 1995 18955
rect 14289 18921 14323 18955
rect 17233 18921 17267 18955
rect 5457 18853 5491 18887
rect 5825 18853 5859 18887
rect 23397 18853 23431 18887
rect 4261 18785 4295 18819
rect 7849 18785 7883 18819
rect 8677 18785 8711 18819
rect 11713 18785 11747 18819
rect 14933 18785 14967 18819
rect 18337 18785 18371 18819
rect 20361 18785 20395 18819
rect 20637 18785 20671 18819
rect 23029 18785 23063 18819
rect 23213 18785 23247 18819
rect 23857 18785 23891 18819
rect 24041 18785 24075 18819
rect 25237 18785 25271 18819
rect 1869 18717 1903 18751
rect 2145 18717 2179 18751
rect 2881 18717 2915 18751
rect 3525 18717 3559 18751
rect 4721 18717 4755 18751
rect 5641 18717 5675 18751
rect 6009 18717 6043 18751
rect 6653 18717 6687 18751
rect 7297 18717 7331 18751
rect 8401 18717 8435 18751
rect 9137 18717 9171 18751
rect 15485 18717 15519 18751
rect 18061 18717 18095 18751
rect 19625 18717 19659 18751
rect 23765 18717 23799 18751
rect 24961 18717 24995 18751
rect 5365 18649 5399 18683
rect 9413 18649 9447 18683
rect 11989 18649 12023 18683
rect 15761 18649 15795 18683
rect 3341 18581 3375 18615
rect 4537 18581 4571 18615
rect 7113 18581 7147 18615
rect 10885 18581 10919 18615
rect 13461 18581 13495 18615
rect 14657 18581 14691 18615
rect 14749 18581 14783 18615
rect 17693 18581 17727 18615
rect 18153 18581 18187 18615
rect 19441 18581 19475 18615
rect 22109 18581 22143 18615
rect 22569 18581 22603 18615
rect 22937 18581 22971 18615
rect 24593 18581 24627 18615
rect 25053 18581 25087 18615
rect 1869 18377 1903 18411
rect 8033 18377 8067 18411
rect 8401 18377 8435 18411
rect 9137 18377 9171 18411
rect 14289 18377 14323 18411
rect 17233 18377 17267 18411
rect 19533 18377 19567 18411
rect 20821 18377 20855 18411
rect 24593 18377 24627 18411
rect 24961 18377 24995 18411
rect 4721 18309 4755 18343
rect 11161 18309 11195 18343
rect 12173 18309 12207 18343
rect 13001 18309 13035 18343
rect 18245 18309 18279 18343
rect 22017 18309 22051 18343
rect 2053 18241 2087 18275
rect 2145 18241 2179 18275
rect 3525 18241 3559 18275
rect 4169 18241 4203 18275
rect 4997 18241 5031 18275
rect 5365 18241 5399 18275
rect 6009 18241 6043 18275
rect 7297 18241 7331 18275
rect 8225 18241 8259 18275
rect 8585 18241 8619 18275
rect 9413 18241 9447 18275
rect 15577 18241 15611 18275
rect 17325 18241 17359 18275
rect 20913 18241 20947 18275
rect 24133 18241 24167 18275
rect 2421 18173 2455 18207
rect 7941 18173 7975 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 15669 18173 15703 18207
rect 15853 18173 15887 18207
rect 17417 18173 17451 18207
rect 21097 18173 21131 18207
rect 25053 18173 25087 18207
rect 25145 18173 25179 18207
rect 3985 18105 4019 18139
rect 4813 18105 4847 18139
rect 5181 18105 5215 18139
rect 5825 18105 5859 18139
rect 16865 18105 16899 18139
rect 23949 18105 23983 18139
rect 7113 18037 7147 18071
rect 11805 18037 11839 18071
rect 15209 18037 15243 18071
rect 20453 18037 20487 18071
rect 23305 18037 23339 18071
rect 2145 17833 2179 17867
rect 5181 17833 5215 17867
rect 6745 17833 6779 17867
rect 7757 17833 7791 17867
rect 8401 17833 8435 17867
rect 16589 17833 16623 17867
rect 18245 17833 18279 17867
rect 7113 17765 7147 17799
rect 9137 17765 9171 17799
rect 11529 17765 11563 17799
rect 13737 17765 13771 17799
rect 11989 17697 12023 17731
rect 12265 17697 12299 17731
rect 14841 17697 14875 17731
rect 17601 17697 17635 17731
rect 19993 17697 20027 17731
rect 20545 17697 20579 17731
rect 22293 17697 22327 17731
rect 23857 17697 23891 17731
rect 2789 17629 2823 17663
rect 3433 17629 3467 17663
rect 4721 17629 4755 17663
rect 6929 17629 6963 17663
rect 7297 17629 7331 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9321 17629 9355 17663
rect 9781 17629 9815 17663
rect 18429 17629 18463 17663
rect 19901 17629 19935 17663
rect 23673 17629 23707 17663
rect 23765 17629 23799 17663
rect 6653 17561 6687 17595
rect 10057 17561 10091 17595
rect 15117 17561 15151 17595
rect 20821 17561 20855 17595
rect 24777 17561 24811 17595
rect 24961 17561 24995 17595
rect 3249 17493 3283 17527
rect 4537 17493 4571 17527
rect 17049 17493 17083 17527
rect 17417 17493 17451 17527
rect 17509 17493 17543 17527
rect 19441 17493 19475 17527
rect 19809 17493 19843 17527
rect 22753 17493 22787 17527
rect 23305 17493 23339 17527
rect 25421 17493 25455 17527
rect 5917 17289 5951 17323
rect 7205 17289 7239 17323
rect 8309 17289 8343 17323
rect 8677 17289 8711 17323
rect 11069 17289 11103 17323
rect 12173 17289 12207 17323
rect 13829 17289 13863 17323
rect 17233 17289 17267 17323
rect 17325 17289 17359 17323
rect 20177 17289 20211 17323
rect 23857 17289 23891 17323
rect 5825 17221 5859 17255
rect 13737 17221 13771 17255
rect 3433 17153 3467 17187
rect 4077 17153 4111 17187
rect 6101 17153 6135 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 8493 17153 8527 17187
rect 8861 17153 8895 17187
rect 9321 17153 9355 17187
rect 12081 17153 12115 17187
rect 14657 17153 14691 17187
rect 15945 17153 15979 17187
rect 18429 17153 18463 17187
rect 20829 17157 20863 17191
rect 21465 17153 21499 17187
rect 22017 17153 22051 17187
rect 22109 17153 22143 17187
rect 24961 17153 24995 17187
rect 8217 17085 8251 17119
rect 9597 17085 9631 17119
rect 12265 17085 12299 17119
rect 13921 17085 13955 17119
rect 16037 17085 16071 17119
rect 16221 17085 16255 17119
rect 17417 17085 17451 17119
rect 18705 17085 18739 17119
rect 22385 17085 22419 17119
rect 3893 17017 3927 17051
rect 14841 17017 14875 17051
rect 15577 17017 15611 17051
rect 25145 17017 25179 17051
rect 4905 16949 4939 16983
rect 6561 16949 6595 16983
rect 11713 16949 11747 16983
rect 13369 16949 13403 16983
rect 16865 16949 16899 16983
rect 20637 16949 20671 16983
rect 21281 16949 21315 16983
rect 21833 16949 21867 16983
rect 24317 16949 24351 16983
rect 4905 16745 4939 16779
rect 10701 16745 10735 16779
rect 11069 16745 11103 16779
rect 16037 16745 16071 16779
rect 16681 16745 16715 16779
rect 19704 16745 19738 16779
rect 21189 16745 21223 16779
rect 6745 16677 6779 16711
rect 7389 16609 7423 16643
rect 7941 16609 7975 16643
rect 11529 16609 11563 16643
rect 12265 16609 12299 16643
rect 14289 16609 14323 16643
rect 14565 16609 14599 16643
rect 17141 16609 17175 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 24869 16609 24903 16643
rect 5641 16541 5675 16575
rect 6285 16541 6319 16575
rect 8585 16541 8619 16575
rect 9597 16541 9631 16575
rect 10241 16541 10275 16575
rect 11989 16541 12023 16575
rect 21833 16541 21867 16575
rect 24685 16473 24719 16507
rect 6101 16405 6135 16439
rect 8401 16405 8435 16439
rect 9413 16405 9447 16439
rect 10057 16405 10091 16439
rect 13737 16405 13771 16439
rect 18889 16405 18923 16439
rect 24041 16405 24075 16439
rect 9137 16201 9171 16235
rect 10609 16201 10643 16235
rect 10977 16201 11011 16235
rect 13461 16201 13495 16235
rect 18521 16201 18555 16235
rect 19441 16201 19475 16235
rect 19901 16201 19935 16235
rect 21097 16201 21131 16235
rect 22477 16201 22511 16235
rect 23857 16201 23891 16235
rect 11989 16133 12023 16167
rect 14381 16133 14415 16167
rect 21189 16133 21223 16167
rect 5181 16065 5215 16099
rect 8493 16065 8527 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 14289 16065 14323 16099
rect 15945 16065 15979 16099
rect 17233 16065 17267 16099
rect 19809 16065 19843 16099
rect 22385 16065 22419 16099
rect 23765 16065 23799 16099
rect 24685 16065 24719 16099
rect 5457 15997 5491 16031
rect 9045 15997 9079 16031
rect 10425 15997 10459 16031
rect 11069 15997 11103 16031
rect 11253 15997 11287 16031
rect 11713 15997 11747 16031
rect 14565 15997 14599 16031
rect 16037 15997 16071 16031
rect 16129 15997 16163 16031
rect 20085 15997 20119 16031
rect 21281 15997 21315 16031
rect 22569 15997 22603 16031
rect 23949 15997 23983 16031
rect 15577 15929 15611 15963
rect 24869 15929 24903 15963
rect 13921 15861 13955 15895
rect 20729 15861 20763 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 16037 15657 16071 15691
rect 18797 15657 18831 15691
rect 20729 15657 20763 15691
rect 9505 15589 9539 15623
rect 12725 15589 12759 15623
rect 19533 15589 19567 15623
rect 9413 15521 9447 15555
rect 10977 15521 11011 15555
rect 13369 15521 13403 15555
rect 14565 15521 14599 15555
rect 17325 15521 17359 15555
rect 20177 15521 20211 15555
rect 21189 15521 21223 15555
rect 21281 15521 21315 15555
rect 24777 15521 24811 15555
rect 9689 15453 9723 15487
rect 10241 15453 10275 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 14289 15453 14323 15487
rect 17049 15453 17083 15487
rect 19901 15453 19935 15487
rect 21097 15453 21131 15487
rect 22201 15453 22235 15487
rect 23581 15453 23615 15487
rect 13093 15385 13127 15419
rect 19993 15385 20027 15419
rect 22017 15385 22051 15419
rect 22753 15385 22787 15419
rect 10333 15317 10367 15351
rect 12449 15317 12483 15351
rect 13185 15317 13219 15351
rect 22845 15317 22879 15351
rect 23397 15317 23431 15351
rect 10977 15113 11011 15147
rect 13461 15113 13495 15147
rect 14841 15113 14875 15147
rect 15485 15113 15519 15147
rect 21189 15113 21223 15147
rect 24685 15113 24719 15147
rect 25145 15113 25179 15147
rect 10517 15045 10551 15079
rect 22109 15045 22143 15079
rect 9873 14977 9907 15011
rect 10793 14977 10827 15011
rect 11161 14977 11195 15011
rect 14105 14977 14139 15011
rect 15025 14977 15059 15011
rect 15669 14977 15703 15011
rect 16313 14977 16347 15011
rect 16865 14977 16899 15011
rect 19441 14977 19475 15011
rect 25329 14977 25363 15011
rect 11713 14909 11747 14943
rect 11989 14909 12023 14943
rect 17141 14909 17175 14943
rect 19717 14909 19751 14943
rect 22937 14909 22971 14943
rect 23213 14909 23247 14943
rect 22293 14841 22327 14875
rect 10609 14773 10643 14807
rect 16129 14773 16163 14807
rect 18613 14773 18647 14807
rect 12449 14569 12483 14603
rect 12909 14569 12943 14603
rect 13277 14569 13311 14603
rect 16037 14501 16071 14535
rect 18245 14501 18279 14535
rect 19441 14501 19475 14535
rect 23305 14501 23339 14535
rect 10977 14433 11011 14467
rect 14289 14433 14323 14467
rect 16773 14433 16807 14467
rect 19993 14433 20027 14467
rect 23949 14433 23983 14467
rect 10701 14365 10735 14399
rect 16497 14365 16531 14399
rect 18889 14365 18923 14399
rect 19809 14365 19843 14399
rect 23673 14365 23707 14399
rect 14565 14297 14599 14331
rect 20821 14297 20855 14331
rect 23765 14297 23799 14331
rect 24685 14297 24719 14331
rect 19901 14229 19935 14263
rect 22109 14229 22143 14263
rect 24777 14229 24811 14263
rect 12725 14025 12759 14059
rect 13185 14025 13219 14059
rect 15761 14025 15795 14059
rect 16129 14025 16163 14059
rect 17049 14025 17083 14059
rect 17509 14025 17543 14059
rect 19533 14025 19567 14059
rect 20729 14025 20763 14059
rect 21097 14025 21131 14059
rect 25237 14025 25271 14059
rect 12265 13957 12299 13991
rect 13829 13957 13863 13991
rect 18245 13957 18279 13991
rect 21189 13957 21223 13991
rect 12541 13889 12575 13923
rect 12909 13889 12943 13923
rect 13369 13889 13403 13923
rect 14013 13889 14047 13923
rect 16313 13889 16347 13923
rect 17417 13889 17451 13923
rect 22017 13889 22051 13923
rect 25145 13889 25179 13923
rect 17693 13821 17727 13855
rect 21281 13821 21315 13855
rect 22293 13821 22327 13855
rect 24041 13821 24075 13855
rect 24501 13821 24535 13855
rect 12357 13753 12391 13787
rect 14276 13685 14310 13719
rect 22109 13685 22143 13719
rect 22556 13685 22590 13719
rect 13553 13481 13587 13515
rect 18245 13481 18279 13515
rect 18889 13481 18923 13515
rect 21465 13481 21499 13515
rect 16037 13413 16071 13447
rect 24593 13413 24627 13447
rect 12081 13345 12115 13379
rect 14289 13345 14323 13379
rect 19717 13345 19751 13379
rect 19993 13345 20027 13379
rect 25053 13345 25087 13379
rect 25145 13345 25179 13379
rect 9597 13277 9631 13311
rect 11805 13277 11839 13311
rect 21925 13277 21959 13311
rect 14565 13209 14599 13243
rect 22201 13209 22235 13243
rect 24961 13209 24995 13243
rect 10885 13141 10919 13175
rect 23673 13141 23707 13175
rect 14657 12937 14691 12971
rect 20821 12937 20855 12971
rect 23765 12937 23799 12971
rect 13185 12869 13219 12903
rect 16681 12869 16715 12903
rect 18797 12869 18831 12903
rect 12909 12801 12943 12835
rect 15117 12801 15151 12835
rect 18521 12801 18555 12835
rect 20729 12801 20763 12835
rect 25053 12801 25087 12835
rect 15393 12733 15427 12767
rect 20913 12733 20947 12767
rect 22017 12733 22051 12767
rect 22293 12733 22327 12767
rect 24409 12733 24443 12767
rect 20269 12665 20303 12699
rect 17969 12597 18003 12631
rect 20361 12597 20395 12631
rect 18153 12393 18187 12427
rect 19704 12393 19738 12427
rect 24041 12393 24075 12427
rect 24777 12393 24811 12427
rect 17509 12325 17543 12359
rect 15761 12257 15795 12291
rect 21833 12257 21867 12291
rect 22569 12257 22603 12291
rect 14289 12189 14323 12223
rect 14565 12189 14599 12223
rect 19441 12189 19475 12223
rect 22293 12189 22327 12223
rect 16037 12121 16071 12155
rect 18705 12121 18739 12155
rect 18889 12121 18923 12155
rect 21741 12121 21775 12155
rect 21189 12053 21223 12087
rect 21281 12053 21315 12087
rect 21649 12053 21683 12087
rect 14473 11849 14507 11883
rect 15117 11849 15151 11883
rect 15853 11849 15887 11883
rect 16129 11849 16163 11883
rect 19165 11849 19199 11883
rect 14013 11781 14047 11815
rect 17141 11781 17175 11815
rect 19625 11781 19659 11815
rect 23305 11781 23339 11815
rect 14657 11713 14691 11747
rect 15301 11713 15335 11747
rect 16313 11713 16347 11747
rect 16865 11713 16899 11747
rect 19349 11713 19383 11747
rect 22017 11713 22051 11747
rect 22109 11713 22143 11747
rect 23949 11713 23983 11747
rect 21097 11645 21131 11679
rect 24777 11645 24811 11679
rect 18613 11509 18647 11543
rect 16497 11305 16531 11339
rect 21833 11305 21867 11339
rect 24593 11305 24627 11339
rect 18889 11237 18923 11271
rect 21189 11237 21223 11271
rect 17141 11169 17175 11203
rect 23857 11169 23891 11203
rect 16037 11101 16071 11135
rect 16681 11101 16715 11135
rect 19993 11101 20027 11135
rect 21373 11101 21407 11135
rect 22017 11101 22051 11135
rect 22661 11101 22695 11135
rect 24777 11101 24811 11135
rect 17417 11033 17451 11067
rect 20177 11033 20211 11067
rect 17325 10761 17359 10795
rect 17693 10761 17727 10795
rect 17233 10693 17267 10727
rect 23305 10693 23339 10727
rect 15209 10625 15243 10659
rect 17509 10625 17543 10659
rect 17877 10625 17911 10659
rect 18613 10625 18647 10659
rect 18981 10625 19015 10659
rect 19625 10625 19659 10659
rect 20269 10625 20303 10659
rect 20913 10625 20947 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 15485 10557 15519 10591
rect 24685 10557 24719 10591
rect 19441 10421 19475 10455
rect 20085 10421 20119 10455
rect 20729 10421 20763 10455
rect 17325 10217 17359 10251
rect 17417 10217 17451 10251
rect 19441 10217 19475 10251
rect 20085 10217 20119 10251
rect 23857 10217 23891 10251
rect 24593 10149 24627 10183
rect 18061 10081 18095 10115
rect 21281 10081 21315 10115
rect 21557 10081 21591 10115
rect 25145 10081 25179 10115
rect 17601 10013 17635 10047
rect 18337 10013 18371 10047
rect 19625 10013 19659 10047
rect 20453 10013 20487 10047
rect 24041 10013 24075 10047
rect 24961 10013 24995 10047
rect 20269 9877 20303 9911
rect 23029 9877 23063 9911
rect 25053 9877 25087 9911
rect 20637 9673 20671 9707
rect 23305 9605 23339 9639
rect 17601 9537 17635 9571
rect 18245 9537 18279 9571
rect 18889 9537 18923 9571
rect 19533 9537 19567 9571
rect 20177 9537 20211 9571
rect 20821 9537 20855 9571
rect 21465 9537 21499 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 24777 9469 24811 9503
rect 19349 9401 19383 9435
rect 19993 9401 20027 9435
rect 18061 9333 18095 9367
rect 18705 9333 18739 9367
rect 21281 9333 21315 9367
rect 11897 9129 11931 9163
rect 21373 9061 21407 9095
rect 10149 8993 10183 9027
rect 19441 8993 19475 9027
rect 23857 8993 23891 9027
rect 19717 8925 19751 8959
rect 20913 8925 20947 8959
rect 21557 8925 21591 8959
rect 22201 8925 22235 8959
rect 22661 8925 22695 8959
rect 10425 8857 10459 8891
rect 24685 8857 24719 8891
rect 24869 8857 24903 8891
rect 20729 8789 20763 8823
rect 22017 8789 22051 8823
rect 19993 8585 20027 8619
rect 21281 8585 21315 8619
rect 23305 8517 23339 8551
rect 20177 8449 20211 8483
rect 20821 8449 20855 8483
rect 21465 8449 21499 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 24593 8381 24627 8415
rect 20637 8313 20671 8347
rect 20729 8041 20763 8075
rect 24593 8041 24627 8075
rect 21373 7973 21407 8007
rect 22201 7973 22235 8007
rect 23857 7905 23891 7939
rect 20913 7837 20947 7871
rect 21557 7837 21591 7871
rect 22845 7837 22879 7871
rect 24777 7837 24811 7871
rect 23305 7429 23339 7463
rect 21465 7361 21499 7395
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 24685 7293 24719 7327
rect 20821 7225 20855 7259
rect 21281 7157 21315 7191
rect 21373 6885 21407 6919
rect 23857 6817 23891 6851
rect 21557 6749 21591 6783
rect 22201 6749 22235 6783
rect 22661 6749 22695 6783
rect 24685 6749 24719 6783
rect 24869 6681 24903 6715
rect 22017 6613 22051 6647
rect 23305 6341 23339 6375
rect 22293 6273 22327 6307
rect 24133 6273 24167 6307
rect 24777 6205 24811 6239
rect 22017 5797 22051 5831
rect 22201 5661 22235 5695
rect 22845 5661 22879 5695
rect 24869 5661 24903 5695
rect 23857 5593 23891 5627
rect 24685 5525 24719 5559
rect 23305 5253 23339 5287
rect 22109 5185 22143 5219
rect 23949 5185 23983 5219
rect 24685 5117 24719 5151
rect 22661 4573 22695 4607
rect 24869 4573 24903 4607
rect 23857 4505 23891 4539
rect 24685 4437 24719 4471
rect 20269 4097 20303 4131
rect 22293 4097 22327 4131
rect 23949 4097 23983 4131
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 24869 3485 24903 3519
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 24685 3349 24719 3383
rect 23305 3077 23339 3111
rect 25145 3077 25179 3111
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 22293 3009 22327 3043
rect 23949 3009 23983 3043
rect 19441 2941 19475 2975
rect 21281 2941 21315 2975
rect 6837 2601 6871 2635
rect 21281 2465 21315 2499
rect 7021 2397 7055 2431
rect 20085 2397 20119 2431
rect 22845 2397 22879 2431
rect 24777 2397 24811 2431
rect 23857 2329 23891 2363
rect 24593 2261 24627 2295
<< metal1 >>
rect 3050 26392 3056 26444
rect 3108 26432 3114 26444
rect 3326 26432 3332 26444
rect 3108 26404 3332 26432
rect 3108 26392 3114 26404
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 2222 26324 2228 26376
rect 2280 26364 2286 26376
rect 22186 26364 22192 26376
rect 2280 26336 22192 26364
rect 2280 26324 2286 26336
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 21450 26296 21456 26308
rect 5276 26268 21456 26296
rect 5276 26240 5304 26268
rect 21450 26256 21456 26268
rect 21508 26256 21514 26308
rect 5258 26188 5264 26240
rect 5316 26188 5322 26240
rect 10226 24896 10232 24948
rect 10284 24936 10290 24948
rect 20714 24936 20720 24948
rect 10284 24908 20720 24936
rect 10284 24896 10290 24908
rect 20714 24896 20720 24908
rect 20772 24896 20778 24948
rect 18506 24828 18512 24880
rect 18564 24868 18570 24880
rect 18782 24868 18788 24880
rect 18564 24840 18788 24868
rect 18564 24828 18570 24840
rect 18782 24828 18788 24840
rect 18840 24828 18846 24880
rect 11514 24760 11520 24812
rect 11572 24800 11578 24812
rect 13446 24800 13452 24812
rect 11572 24772 13452 24800
rect 11572 24760 11578 24772
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 23382 24800 23388 24812
rect 14240 24772 23388 24800
rect 14240 24760 14246 24772
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 6546 24692 6552 24744
rect 6604 24732 6610 24744
rect 13906 24732 13912 24744
rect 6604 24704 13912 24732
rect 6604 24692 6610 24704
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 16574 24692 16580 24744
rect 16632 24732 16638 24744
rect 21082 24732 21088 24744
rect 16632 24704 21088 24732
rect 16632 24692 16638 24704
rect 21082 24692 21088 24704
rect 21140 24692 21146 24744
rect 4890 24624 4896 24676
rect 4948 24664 4954 24676
rect 14734 24664 14740 24676
rect 4948 24636 14740 24664
rect 4948 24624 4954 24636
rect 14734 24624 14740 24636
rect 14792 24624 14798 24676
rect 16022 24624 16028 24676
rect 16080 24664 16086 24676
rect 22002 24664 22008 24676
rect 16080 24636 22008 24664
rect 16080 24624 16086 24636
rect 22002 24624 22008 24636
rect 22060 24624 22066 24676
rect 4798 24556 4804 24608
rect 4856 24596 4862 24608
rect 15470 24596 15476 24608
rect 4856 24568 15476 24596
rect 4856 24556 4862 24568
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 16390 24556 16396 24608
rect 16448 24596 16454 24608
rect 24210 24596 24216 24608
rect 16448 24568 24216 24596
rect 16448 24556 16454 24568
rect 24210 24556 24216 24568
rect 24268 24556 24274 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 15470 24352 15476 24404
rect 15528 24352 15534 24404
rect 17589 24395 17647 24401
rect 17589 24392 17601 24395
rect 15856 24364 17601 24392
rect 12710 24284 12716 24336
rect 12768 24324 12774 24336
rect 15856 24324 15884 24364
rect 17589 24361 17601 24364
rect 17635 24392 17647 24395
rect 18506 24392 18512 24404
rect 17635 24364 18512 24392
rect 17635 24361 17647 24364
rect 17589 24355 17647 24361
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 21818 24392 21824 24404
rect 20088 24364 21824 24392
rect 18141 24327 18199 24333
rect 18141 24324 18153 24327
rect 12768 24296 15884 24324
rect 15948 24296 18153 24324
rect 12768 24284 12774 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6454 24256 6460 24268
rect 3283 24228 6460 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 8205 24259 8263 24265
rect 6564 24228 7236 24256
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 3878 24188 3884 24200
rect 2271 24160 3884 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 5442 24148 5448 24200
rect 5500 24188 5506 24200
rect 6564 24188 6592 24228
rect 5500 24160 6592 24188
rect 6733 24191 6791 24197
rect 5500 24148 5506 24160
rect 6733 24157 6745 24191
rect 6779 24188 6791 24191
rect 7006 24188 7012 24200
rect 6779 24160 7012 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 7006 24148 7012 24160
rect 7064 24148 7070 24200
rect 7208 24197 7236 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9674 24256 9680 24268
rect 8251 24228 9680 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10962 24216 10968 24268
rect 11020 24216 11026 24268
rect 12434 24216 12440 24268
rect 12492 24256 12498 24268
rect 12805 24259 12863 24265
rect 12805 24256 12817 24259
rect 12492 24228 12817 24256
rect 12492 24216 12498 24228
rect 12805 24225 12817 24228
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 13906 24216 13912 24268
rect 13964 24256 13970 24268
rect 15948 24256 15976 24296
rect 18141 24293 18153 24296
rect 18187 24293 18199 24327
rect 19794 24324 19800 24336
rect 18141 24287 18199 24293
rect 18432 24296 19800 24324
rect 13964 24228 15976 24256
rect 13964 24216 13970 24228
rect 16114 24216 16120 24268
rect 16172 24256 16178 24268
rect 16209 24259 16267 24265
rect 16209 24256 16221 24259
rect 16172 24228 16221 24256
rect 16172 24216 16178 24228
rect 16209 24225 16221 24228
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 16390 24216 16396 24268
rect 16448 24216 16454 24268
rect 18432 24256 18460 24296
rect 19794 24284 19800 24296
rect 19852 24284 19858 24336
rect 17420 24228 18460 24256
rect 18785 24259 18843 24265
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 8662 24120 8668 24132
rect 5859 24092 8668 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 9324 24120 9352 24151
rect 9582 24148 9588 24200
rect 9640 24188 9646 24200
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 9640 24160 9781 24188
rect 9640 24148 9646 24160
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 11882 24148 11888 24200
rect 11940 24148 11946 24200
rect 12526 24148 12532 24200
rect 12584 24148 12590 24200
rect 13722 24148 13728 24200
rect 13780 24188 13786 24200
rect 16945 24191 17003 24197
rect 16945 24188 16957 24191
rect 13780 24160 16957 24188
rect 13780 24148 13786 24160
rect 16945 24157 16957 24160
rect 16991 24157 17003 24191
rect 16945 24151 17003 24157
rect 14274 24120 14280 24132
rect 9324 24092 14280 24120
rect 14274 24080 14280 24092
rect 14332 24080 14338 24132
rect 14366 24080 14372 24132
rect 14424 24080 14430 24132
rect 14550 24080 14556 24132
rect 14608 24120 14614 24132
rect 15381 24123 15439 24129
rect 15381 24120 15393 24123
rect 14608 24092 15393 24120
rect 14608 24080 14614 24092
rect 15381 24089 15393 24092
rect 15427 24089 15439 24123
rect 15381 24083 15439 24089
rect 15764 24092 16712 24120
rect 3694 24012 3700 24064
rect 3752 24052 3758 24064
rect 3973 24055 4031 24061
rect 3973 24052 3985 24055
rect 3752 24024 3985 24052
rect 3752 24012 3758 24024
rect 3973 24021 3985 24024
rect 4019 24021 4031 24055
rect 3973 24015 4031 24021
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 7098 24052 7104 24064
rect 6595 24024 7104 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 15764 24061 15792 24092
rect 14461 24055 14519 24061
rect 14461 24052 14473 24055
rect 9732 24024 14473 24052
rect 9732 24012 9738 24024
rect 14461 24021 14473 24024
rect 14507 24021 14519 24055
rect 14461 24015 14519 24021
rect 15749 24055 15807 24061
rect 15749 24021 15761 24055
rect 15795 24021 15807 24055
rect 15749 24015 15807 24021
rect 16117 24055 16175 24061
rect 16117 24021 16129 24055
rect 16163 24052 16175 24055
rect 16574 24052 16580 24064
rect 16163 24024 16580 24052
rect 16163 24021 16175 24024
rect 16117 24015 16175 24021
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 16684 24052 16712 24092
rect 16758 24080 16764 24132
rect 16816 24080 16822 24132
rect 17420 24052 17448 24228
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 19150 24256 19156 24268
rect 18831 24228 19156 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 20088 24265 20116 24364
rect 21818 24352 21824 24364
rect 21876 24352 21882 24404
rect 20714 24284 20720 24336
rect 20772 24324 20778 24336
rect 23753 24327 23811 24333
rect 23753 24324 23765 24327
rect 20772 24296 23765 24324
rect 20772 24284 20778 24296
rect 23753 24293 23765 24296
rect 23799 24324 23811 24327
rect 23799 24296 24992 24324
rect 23799 24293 23811 24296
rect 23753 24287 23811 24293
rect 20073 24259 20131 24265
rect 20073 24225 20085 24259
rect 20119 24225 20131 24259
rect 20073 24219 20131 24225
rect 20809 24259 20867 24265
rect 20809 24225 20821 24259
rect 20855 24256 20867 24259
rect 21910 24256 21916 24268
rect 20855 24228 21916 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 21910 24216 21916 24228
rect 21968 24216 21974 24268
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24188 19855 24191
rect 20438 24188 20444 24200
rect 19843 24160 20444 24188
rect 19843 24157 19855 24160
rect 19797 24151 19855 24157
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 21082 24148 21088 24200
rect 21140 24188 21146 24200
rect 21358 24188 21364 24200
rect 21140 24160 21364 24188
rect 21140 24148 21146 24160
rect 21358 24148 21364 24160
rect 21416 24148 21422 24200
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24188 22063 24191
rect 24486 24188 24492 24200
rect 22051 24160 24492 24188
rect 22051 24157 22063 24160
rect 22005 24151 22063 24157
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 24964 24197 24992 24296
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 24949 24191 25007 24197
rect 24949 24157 24961 24191
rect 24995 24157 25007 24191
rect 24949 24151 25007 24157
rect 17494 24080 17500 24132
rect 17552 24120 17558 24132
rect 22554 24120 22560 24132
rect 17552 24092 22560 24120
rect 17552 24080 17558 24092
rect 22554 24080 22560 24092
rect 22612 24080 22618 24132
rect 22830 24080 22836 24132
rect 22888 24080 22894 24132
rect 23842 24080 23848 24132
rect 23900 24120 23906 24132
rect 25148 24120 25176 24219
rect 23900 24092 25176 24120
rect 23900 24080 23906 24092
rect 16684 24024 17448 24052
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 19334 24052 19340 24064
rect 18647 24024 19340 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 19334 24012 19340 24024
rect 19392 24012 19398 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 20625 24055 20683 24061
rect 20625 24052 20637 24055
rect 19944 24024 20637 24052
rect 19944 24012 19950 24024
rect 20625 24021 20637 24024
rect 20671 24021 20683 24055
rect 20625 24015 20683 24021
rect 23934 24012 23940 24064
rect 23992 24052 23998 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 23992 24024 24593 24052
rect 23992 24012 23998 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 25038 24012 25044 24064
rect 25096 24012 25102 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 4212 23820 11836 23848
rect 4212 23808 4218 23820
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 5074 23780 5080 23792
rect 4019 23752 5080 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 5074 23740 5080 23752
rect 5132 23740 5138 23792
rect 5813 23783 5871 23789
rect 5813 23749 5825 23783
rect 5859 23780 5871 23783
rect 7558 23780 7564 23792
rect 5859 23752 7564 23780
rect 5859 23749 5871 23752
rect 5813 23743 5871 23749
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 10134 23780 10140 23792
rect 9171 23752 10140 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 10134 23740 10140 23752
rect 10192 23740 10198 23792
rect 10870 23740 10876 23792
rect 10928 23740 10934 23792
rect 11808 23780 11836 23820
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 14274 23848 14280 23860
rect 11940 23820 14280 23848
rect 11940 23808 11946 23820
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 16853 23851 16911 23857
rect 16853 23817 16865 23851
rect 16899 23848 16911 23851
rect 25038 23848 25044 23860
rect 16899 23820 25044 23848
rect 16899 23817 16911 23820
rect 16853 23811 16911 23817
rect 25038 23808 25044 23820
rect 25096 23808 25102 23860
rect 14461 23783 14519 23789
rect 11808 23752 12204 23780
rect 934 23672 940 23724
rect 992 23712 998 23724
rect 1673 23715 1731 23721
rect 1673 23712 1685 23715
rect 992 23684 1685 23712
rect 992 23672 998 23684
rect 1673 23681 1685 23684
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 4890 23712 4896 23724
rect 4847 23684 4896 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 2976 23644 3004 23675
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 6546 23672 6552 23724
rect 6604 23672 6610 23724
rect 6656 23684 7236 23712
rect 6656 23644 6684 23684
rect 2976 23616 6684 23644
rect 6730 23604 6736 23656
rect 6788 23644 6794 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6788 23616 6837 23644
rect 6788 23604 6794 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 7208 23644 7236 23684
rect 7282 23672 7288 23724
rect 7340 23712 7346 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7340 23684 7941 23712
rect 7340 23672 7346 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 8386 23672 8392 23724
rect 8444 23712 8450 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 8444 23684 9781 23712
rect 8444 23672 8450 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 9769 23675 9827 23681
rect 9876 23684 12081 23712
rect 8478 23644 8484 23656
rect 7208 23616 8484 23644
rect 6825 23607 6883 23613
rect 8478 23604 8484 23616
rect 8536 23604 8542 23656
rect 4338 23536 4344 23588
rect 4396 23576 4402 23588
rect 9876 23576 9904 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 4396 23548 9904 23576
rect 12176 23576 12204 23752
rect 14461 23749 14473 23783
rect 14507 23780 14519 23783
rect 17126 23780 17132 23792
rect 14507 23752 17132 23780
rect 14507 23749 14519 23752
rect 14461 23743 14519 23749
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 17221 23783 17279 23789
rect 17221 23749 17233 23783
rect 17267 23780 17279 23783
rect 18414 23780 18420 23792
rect 17267 23752 18420 23780
rect 17267 23749 17279 23752
rect 17221 23743 17279 23749
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 18690 23740 18696 23792
rect 18748 23740 18754 23792
rect 22462 23780 22468 23792
rect 20640 23752 22468 23780
rect 14274 23672 14280 23724
rect 14332 23712 14338 23724
rect 20640 23721 20668 23752
rect 22462 23740 22468 23752
rect 22520 23740 22526 23792
rect 22830 23740 22836 23792
rect 22888 23740 22894 23792
rect 24762 23740 24768 23792
rect 24820 23780 24826 23792
rect 25133 23783 25191 23789
rect 25133 23780 25145 23783
rect 24820 23752 25145 23780
rect 24820 23740 24826 23752
rect 25133 23749 25145 23752
rect 25179 23749 25191 23783
rect 25133 23743 25191 23749
rect 14369 23715 14427 23721
rect 14369 23712 14381 23715
rect 14332 23684 14381 23712
rect 14332 23672 14338 23684
rect 14369 23681 14381 23684
rect 14415 23681 14427 23715
rect 14369 23675 14427 23681
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 20165 23715 20223 23721
rect 20165 23681 20177 23715
rect 20211 23712 20223 23715
rect 20625 23715 20683 23721
rect 20625 23712 20637 23715
rect 20211 23684 20637 23712
rect 20211 23681 20223 23684
rect 20165 23675 20223 23681
rect 20625 23681 20637 23684
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 12250 23604 12256 23656
rect 12308 23644 12314 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12308 23616 12541 23644
rect 12308 23604 12314 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 14550 23604 14556 23656
rect 14608 23604 14614 23656
rect 14001 23579 14059 23585
rect 14001 23576 14013 23579
rect 12176 23548 14013 23576
rect 4396 23536 4402 23548
rect 14001 23545 14013 23548
rect 14047 23545 14059 23579
rect 14001 23539 14059 23545
rect 15565 23579 15623 23585
rect 15565 23545 15577 23579
rect 15611 23545 15623 23579
rect 15565 23539 15623 23545
rect 1765 23511 1823 23517
rect 1765 23477 1777 23511
rect 1811 23508 1823 23511
rect 6546 23508 6552 23520
rect 1811 23480 6552 23508
rect 1811 23477 1823 23480
rect 1765 23471 1823 23477
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 7006 23468 7012 23520
rect 7064 23508 7070 23520
rect 15580 23508 15608 23539
rect 7064 23480 15608 23508
rect 15948 23508 15976 23675
rect 22002 23672 22008 23724
rect 22060 23672 22066 23724
rect 16022 23604 16028 23656
rect 16080 23604 16086 23656
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 16209 23647 16267 23653
rect 16209 23644 16221 23647
rect 16172 23616 16221 23644
rect 16172 23604 16178 23616
rect 16209 23613 16221 23616
rect 16255 23644 16267 23647
rect 16298 23644 16304 23656
rect 16255 23616 16304 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 16298 23604 16304 23616
rect 16356 23604 16362 23656
rect 17310 23604 17316 23656
rect 17368 23604 17374 23656
rect 17494 23604 17500 23656
rect 17552 23604 17558 23656
rect 17862 23604 17868 23656
rect 17920 23604 17926 23656
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23644 18199 23647
rect 19150 23644 19156 23656
rect 18187 23616 19156 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 19150 23604 19156 23616
rect 19208 23604 19214 23656
rect 20901 23647 20959 23653
rect 20901 23644 20913 23647
rect 19260 23616 20913 23644
rect 19260 23588 19288 23616
rect 20901 23613 20913 23616
rect 20947 23644 20959 23647
rect 21266 23644 21272 23656
rect 20947 23616 21272 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 21266 23604 21272 23616
rect 21324 23604 21330 23656
rect 22094 23604 22100 23656
rect 22152 23604 22158 23656
rect 22373 23647 22431 23653
rect 22373 23613 22385 23647
rect 22419 23644 22431 23647
rect 22462 23644 22468 23656
rect 22419 23616 22468 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 23842 23604 23848 23656
rect 23900 23604 23906 23656
rect 19242 23536 19248 23588
rect 19300 23536 19306 23588
rect 19702 23536 19708 23588
rect 19760 23576 19766 23588
rect 20162 23576 20168 23588
rect 19760 23548 20168 23576
rect 19760 23536 19766 23548
rect 20162 23536 20168 23548
rect 20220 23536 20226 23588
rect 25590 23576 25596 23588
rect 23860 23548 25596 23576
rect 18874 23508 18880 23520
rect 15948 23480 18880 23508
rect 7064 23468 7070 23480
rect 18874 23468 18880 23480
rect 18932 23468 18938 23520
rect 19610 23468 19616 23520
rect 19668 23468 19674 23520
rect 19794 23468 19800 23520
rect 19852 23508 19858 23520
rect 20346 23508 20352 23520
rect 19852 23480 20352 23508
rect 19852 23468 19858 23480
rect 20346 23468 20352 23480
rect 20404 23468 20410 23520
rect 21821 23511 21879 23517
rect 21821 23477 21833 23511
rect 21867 23508 21879 23511
rect 23860 23508 23888 23548
rect 25590 23536 25596 23548
rect 25648 23536 25654 23588
rect 21867 23480 23888 23508
rect 21867 23477 21879 23480
rect 21821 23471 21879 23477
rect 25222 23468 25228 23520
rect 25280 23468 25286 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 9674 23304 9680 23316
rect 4212 23276 9680 23304
rect 4212 23264 4218 23276
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 9950 23264 9956 23316
rect 10008 23304 10014 23316
rect 14918 23304 14924 23316
rect 10008 23276 14924 23304
rect 10008 23264 10014 23276
rect 14918 23264 14924 23276
rect 14976 23264 14982 23316
rect 16298 23264 16304 23316
rect 16356 23304 16362 23316
rect 18877 23307 18935 23313
rect 18877 23304 18889 23307
rect 16356 23276 18889 23304
rect 16356 23264 16362 23276
rect 18877 23273 18889 23276
rect 18923 23273 18935 23307
rect 18877 23267 18935 23273
rect 19150 23264 19156 23316
rect 19208 23304 19214 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 19208 23276 21189 23304
rect 19208 23264 19214 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 22002 23304 22008 23316
rect 21177 23267 21235 23273
rect 21560 23276 22008 23304
rect 5074 23196 5080 23248
rect 5132 23236 5138 23248
rect 5350 23236 5356 23248
rect 5132 23208 5356 23236
rect 5132 23196 5138 23208
rect 5350 23196 5356 23208
rect 5408 23196 5414 23248
rect 7650 23236 7656 23248
rect 6564 23208 7656 23236
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 4614 23168 4620 23180
rect 3283 23140 4620 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 6564 23177 6592 23208
rect 7650 23196 7656 23208
rect 7708 23196 7714 23248
rect 9398 23236 9404 23248
rect 8220 23208 9404 23236
rect 6549 23171 6607 23177
rect 5368 23140 6500 23168
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 3602 23100 3608 23112
rect 2271 23072 3608 23100
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 3602 23060 3608 23072
rect 3660 23060 3666 23112
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4338 23100 4344 23112
rect 4295 23072 4344 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 3988 23032 4016 23063
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 5368 23032 5396 23140
rect 5537 23103 5595 23109
rect 5537 23069 5549 23103
rect 5583 23100 5595 23103
rect 5626 23100 5632 23112
rect 5583 23072 5632 23100
rect 5583 23069 5595 23072
rect 5537 23063 5595 23069
rect 5626 23060 5632 23072
rect 5684 23060 5690 23112
rect 3988 23004 5396 23032
rect 6472 23032 6500 23140
rect 6549 23137 6561 23171
rect 6595 23137 6607 23171
rect 7374 23168 7380 23180
rect 6549 23131 6607 23137
rect 7208 23140 7380 23168
rect 7208 23109 7236 23140
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 8220 23177 8248 23208
rect 9398 23196 9404 23208
rect 9456 23196 9462 23248
rect 10134 23196 10140 23248
rect 10192 23236 10198 23248
rect 13906 23236 13912 23248
rect 10192 23208 13912 23236
rect 10192 23196 10198 23208
rect 13906 23196 13912 23208
rect 13964 23196 13970 23248
rect 18506 23196 18512 23248
rect 18564 23236 18570 23248
rect 18564 23208 19564 23236
rect 18564 23196 18570 23208
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23137 8263 23171
rect 8205 23131 8263 23137
rect 8570 23128 8576 23180
rect 8628 23168 8634 23180
rect 8628 23140 9904 23168
rect 8628 23128 8634 23140
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23100 9459 23103
rect 9766 23100 9772 23112
rect 9447 23072 9772 23100
rect 9447 23069 9459 23072
rect 9401 23063 9459 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 9876 23109 9904 23140
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11664 23140 12173 23168
rect 11664 23128 11670 23140
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 12161 23131 12219 23137
rect 13538 23128 13544 23180
rect 13596 23168 13602 23180
rect 14921 23171 14979 23177
rect 14921 23168 14933 23171
rect 13596 23140 14933 23168
rect 13596 23128 13602 23140
rect 14921 23137 14933 23140
rect 14967 23137 14979 23171
rect 14921 23131 14979 23137
rect 15197 23171 15255 23177
rect 15197 23137 15209 23171
rect 15243 23168 15255 23171
rect 15930 23168 15936 23180
rect 15243 23140 15936 23168
rect 15243 23137 15255 23140
rect 15197 23131 15255 23137
rect 15930 23128 15936 23140
rect 15988 23128 15994 23180
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23168 17187 23171
rect 17862 23168 17868 23180
rect 17175 23140 17868 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 17862 23128 17868 23140
rect 17920 23168 17926 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 17920 23140 19441 23168
rect 17920 23128 17926 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19536 23168 19564 23208
rect 21450 23196 21456 23248
rect 21508 23196 21514 23248
rect 21468 23168 21496 23196
rect 21560 23177 21588 23276
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 22278 23264 22284 23316
rect 22336 23304 22342 23316
rect 24026 23304 24032 23316
rect 22336 23276 24032 23304
rect 22336 23264 22342 23276
rect 24026 23264 24032 23276
rect 24084 23264 24090 23316
rect 23198 23196 23204 23248
rect 23256 23236 23262 23248
rect 24946 23236 24952 23248
rect 23256 23208 24952 23236
rect 23256 23196 23262 23208
rect 24946 23196 24952 23208
rect 25004 23196 25010 23248
rect 19536 23140 21496 23168
rect 21545 23171 21603 23177
rect 19429 23131 19487 23137
rect 21545 23137 21557 23171
rect 21591 23137 21603 23171
rect 21545 23131 21603 23137
rect 21818 23128 21824 23180
rect 21876 23168 21882 23180
rect 22278 23168 22284 23180
rect 21876 23140 22284 23168
rect 21876 23128 21882 23140
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 25133 23171 25191 23177
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 11698 23060 11704 23112
rect 11756 23060 11762 23112
rect 13725 23103 13783 23109
rect 13725 23069 13737 23103
rect 13771 23069 13783 23103
rect 13725 23063 13783 23069
rect 13740 23032 13768 23063
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23069 21511 23103
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 21453 23063 21511 23069
rect 23768 23072 24961 23100
rect 15470 23032 15476 23044
rect 6472 23004 11928 23032
rect 13740 23004 15476 23032
rect 1946 22924 1952 22976
rect 2004 22964 2010 22976
rect 4154 22964 4160 22976
rect 2004 22936 4160 22964
rect 2004 22924 2010 22936
rect 4154 22924 4160 22936
rect 4212 22924 4218 22976
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 11698 22964 11704 22976
rect 9263 22936 11704 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 11900 22964 11928 23004
rect 15470 22992 15476 23004
rect 15528 22992 15534 23044
rect 15654 22992 15660 23044
rect 15712 22992 15718 23044
rect 17412 23035 17470 23041
rect 17412 23001 17424 23035
rect 17458 23001 17470 23035
rect 17412 22995 17470 23001
rect 13541 22967 13599 22973
rect 13541 22964 13553 22967
rect 11900 22936 13553 22964
rect 13541 22933 13553 22936
rect 13587 22933 13599 22967
rect 13541 22927 13599 22933
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 16669 22967 16727 22973
rect 16669 22964 16681 22967
rect 14148 22936 16681 22964
rect 14148 22924 14154 22936
rect 16669 22933 16681 22936
rect 16715 22964 16727 22967
rect 17218 22964 17224 22976
rect 16715 22936 17224 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 17218 22924 17224 22936
rect 17276 22924 17282 22976
rect 17420 22964 17448 22995
rect 17954 22992 17960 23044
rect 18012 22992 18018 23044
rect 19242 22992 19248 23044
rect 19300 23032 19306 23044
rect 19300 23004 19656 23032
rect 19300 22992 19306 23004
rect 19628 22976 19656 23004
rect 19702 22992 19708 23044
rect 19760 22992 19766 23044
rect 19978 22992 19984 23044
rect 20036 23032 20042 23044
rect 20036 23004 20194 23032
rect 20036 22992 20042 23004
rect 17494 22964 17500 22976
rect 17420 22936 17500 22964
rect 17494 22924 17500 22936
rect 17552 22964 17558 22976
rect 19518 22964 19524 22976
rect 17552 22936 19524 22964
rect 17552 22924 17558 22936
rect 19518 22924 19524 22936
rect 19576 22924 19582 22976
rect 19610 22924 19616 22976
rect 19668 22924 19674 22976
rect 21468 22964 21496 23063
rect 21910 22992 21916 23044
rect 21968 23032 21974 23044
rect 21968 23004 22310 23032
rect 21968 22992 21974 23004
rect 21634 22964 21640 22976
rect 21468 22936 21640 22964
rect 21634 22924 21640 22936
rect 21692 22924 21698 22976
rect 21726 22924 21732 22976
rect 21784 22964 21790 22976
rect 22002 22964 22008 22976
rect 21784 22936 22008 22964
rect 21784 22924 21790 22936
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 22204 22964 22232 23004
rect 23106 22992 23112 23044
rect 23164 23032 23170 23044
rect 23768 23041 23796 23072
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 23753 23035 23811 23041
rect 23753 23032 23765 23035
rect 23164 23004 23765 23032
rect 23164 22992 23170 23004
rect 23753 23001 23765 23004
rect 23799 23001 23811 23035
rect 23753 22995 23811 23001
rect 24026 22992 24032 23044
rect 24084 23032 24090 23044
rect 25148 23032 25176 23131
rect 24084 23004 25176 23032
rect 24084 22992 24090 23004
rect 22830 22964 22836 22976
rect 22204 22936 22836 22964
rect 22830 22924 22836 22936
rect 22888 22924 22894 22976
rect 23293 22967 23351 22973
rect 23293 22933 23305 22967
rect 23339 22964 23351 22967
rect 23382 22964 23388 22976
rect 23339 22936 23388 22964
rect 23339 22933 23351 22936
rect 23293 22927 23351 22933
rect 23382 22924 23388 22936
rect 23440 22924 23446 22976
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22964 24639 22967
rect 24854 22964 24860 22976
rect 24627 22936 24860 22964
rect 24627 22933 24639 22936
rect 24581 22927 24639 22933
rect 24854 22924 24860 22936
rect 24912 22924 24918 22976
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25406 22964 25412 22976
rect 25087 22936 25412 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 25406 22924 25412 22936
rect 25464 22924 25470 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 8570 22760 8576 22772
rect 4448 22732 8576 22760
rect 4448 22704 4476 22732
rect 8570 22720 8576 22732
rect 8628 22720 8634 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 9548 22732 11713 22760
rect 9548 22720 9554 22732
rect 11701 22729 11713 22732
rect 11747 22729 11759 22763
rect 11701 22723 11759 22729
rect 12161 22763 12219 22769
rect 12161 22729 12173 22763
rect 12207 22760 12219 22763
rect 12207 22732 13492 22760
rect 12207 22729 12219 22732
rect 12161 22723 12219 22729
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4246 22692 4252 22704
rect 4019 22664 4252 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 4430 22652 4436 22704
rect 4488 22652 4494 22704
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 9950 22692 9956 22704
rect 8864 22664 9956 22692
rect 934 22584 940 22636
rect 992 22624 998 22636
rect 1673 22627 1731 22633
rect 1673 22624 1685 22627
rect 992 22596 1685 22624
rect 992 22584 998 22596
rect 1673 22593 1685 22596
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 4522 22624 4528 22636
rect 3007 22596 4528 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 4522 22584 4528 22596
rect 4580 22584 4586 22636
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22624 4859 22627
rect 5166 22624 5172 22636
rect 4847 22596 5172 22624
rect 4847 22593 4859 22596
rect 4801 22587 4859 22593
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 6638 22584 6644 22636
rect 6696 22584 6702 22636
rect 6822 22584 6828 22636
rect 6880 22624 6886 22636
rect 7561 22627 7619 22633
rect 7561 22624 7573 22627
rect 6880 22596 7573 22624
rect 6880 22584 6886 22596
rect 7561 22593 7573 22596
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 8864 22624 8892 22664
rect 9950 22652 9956 22664
rect 10008 22652 10014 22704
rect 11330 22692 11336 22704
rect 10902 22664 11336 22692
rect 11330 22652 11336 22664
rect 11388 22652 11394 22704
rect 12250 22652 12256 22704
rect 12308 22692 12314 22704
rect 12618 22692 12624 22704
rect 12308 22664 12624 22692
rect 12308 22652 12314 22664
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 7800 22596 8892 22624
rect 7800 22584 7806 22596
rect 11422 22584 11428 22636
rect 11480 22624 11486 22636
rect 12069 22627 12127 22633
rect 12069 22624 12081 22627
rect 11480 22596 12081 22624
rect 11480 22584 11486 22596
rect 12069 22593 12081 22596
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 13081 22627 13139 22633
rect 13081 22593 13093 22627
rect 13127 22624 13139 22627
rect 13354 22624 13360 22636
rect 13127 22596 13360 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9180 22528 9413 22556
rect 9180 22516 9186 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 12158 22556 12164 22568
rect 9723 22528 12164 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 12158 22516 12164 22528
rect 12216 22556 12222 22568
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 12216 22528 12265 22556
rect 12216 22516 12222 22528
rect 12253 22525 12265 22528
rect 12299 22525 12311 22559
rect 12253 22519 12311 22525
rect 12342 22516 12348 22568
rect 12400 22556 12406 22568
rect 13464 22556 13492 22732
rect 14550 22720 14556 22772
rect 14608 22760 14614 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 14608 22732 15301 22760
rect 14608 22720 14614 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 15930 22720 15936 22772
rect 15988 22720 15994 22772
rect 17034 22720 17040 22772
rect 17092 22720 17098 22772
rect 17126 22720 17132 22772
rect 17184 22760 17190 22772
rect 17221 22763 17279 22769
rect 17221 22760 17233 22763
rect 17184 22732 17233 22760
rect 17184 22720 17190 22732
rect 17221 22729 17233 22732
rect 17267 22729 17279 22763
rect 17221 22723 17279 22729
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 18506 22760 18512 22772
rect 17460 22732 18512 22760
rect 17460 22720 17466 22732
rect 18506 22720 18512 22732
rect 18564 22720 18570 22772
rect 18874 22720 18880 22772
rect 18932 22760 18938 22772
rect 18969 22763 19027 22769
rect 18969 22760 18981 22763
rect 18932 22732 18981 22760
rect 18932 22720 18938 22732
rect 18969 22729 18981 22732
rect 19015 22729 19027 22763
rect 18969 22723 19027 22729
rect 19978 22720 19984 22772
rect 20036 22760 20042 22772
rect 20165 22763 20223 22769
rect 20165 22760 20177 22763
rect 20036 22732 20177 22760
rect 20036 22720 20042 22732
rect 20165 22729 20177 22732
rect 20211 22729 20223 22763
rect 20165 22723 20223 22729
rect 22002 22720 22008 22772
rect 22060 22760 22066 22772
rect 22278 22760 22284 22772
rect 22060 22732 22284 22760
rect 22060 22720 22066 22732
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 22373 22763 22431 22769
rect 22373 22729 22385 22763
rect 22419 22760 22431 22763
rect 25222 22760 25228 22772
rect 22419 22732 25228 22760
rect 22419 22729 22431 22732
rect 22373 22723 22431 22729
rect 13817 22695 13875 22701
rect 13817 22661 13829 22695
rect 13863 22692 13875 22695
rect 14090 22692 14096 22704
rect 13863 22664 14096 22692
rect 13863 22661 13875 22664
rect 13817 22655 13875 22661
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 14274 22652 14280 22704
rect 14332 22652 14338 22704
rect 16482 22652 16488 22704
rect 16540 22692 16546 22704
rect 17589 22695 17647 22701
rect 17589 22692 17601 22695
rect 16540 22664 17601 22692
rect 16540 22652 16546 22664
rect 17589 22661 17601 22664
rect 17635 22661 17647 22695
rect 17589 22655 17647 22661
rect 19150 22652 19156 22704
rect 19208 22692 19214 22704
rect 20254 22692 20260 22704
rect 19208 22664 20260 22692
rect 19208 22652 19214 22664
rect 20254 22652 20260 22664
rect 20312 22652 20318 22704
rect 20438 22652 20444 22704
rect 20496 22692 20502 22704
rect 22388 22692 22416 22723
rect 25222 22720 25228 22732
rect 25280 22720 25286 22772
rect 20496 22664 22416 22692
rect 20496 22652 20502 22664
rect 21836 22636 21864 22664
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 15102 22584 15108 22636
rect 15160 22584 15166 22636
rect 15746 22584 15752 22636
rect 15804 22624 15810 22636
rect 15841 22627 15899 22633
rect 15841 22624 15853 22627
rect 15804 22596 15853 22624
rect 15804 22584 15810 22596
rect 15841 22593 15853 22596
rect 15887 22593 15899 22627
rect 16850 22624 16856 22636
rect 15841 22587 15899 22593
rect 15948 22596 16856 22624
rect 15120 22556 15148 22584
rect 12400 22528 13400 22556
rect 13464 22528 15148 22556
rect 12400 22516 12406 22528
rect 1857 22491 1915 22497
rect 1857 22457 1869 22491
rect 1903 22488 1915 22491
rect 7006 22488 7012 22500
rect 1903 22460 7012 22488
rect 1903 22457 1915 22460
rect 1857 22451 1915 22457
rect 7006 22448 7012 22460
rect 7064 22448 7070 22500
rect 11146 22448 11152 22500
rect 11204 22488 11210 22500
rect 11882 22488 11888 22500
rect 11204 22460 11888 22488
rect 11204 22448 11210 22460
rect 11882 22448 11888 22460
rect 11940 22448 11946 22500
rect 6730 22380 6736 22432
rect 6788 22380 6794 22432
rect 9306 22380 9312 22432
rect 9364 22420 9370 22432
rect 12250 22420 12256 22432
rect 9364 22392 12256 22420
rect 9364 22380 9370 22392
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 12618 22380 12624 22432
rect 12676 22420 12682 22432
rect 12897 22423 12955 22429
rect 12897 22420 12909 22423
rect 12676 22392 12909 22420
rect 12676 22380 12682 22392
rect 12897 22389 12909 22392
rect 12943 22389 12955 22423
rect 13372 22420 13400 22528
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 15948 22556 15976 22596
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 16945 22627 17003 22633
rect 16945 22593 16957 22627
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 15620 22528 15976 22556
rect 15620 22516 15626 22528
rect 16298 22516 16304 22568
rect 16356 22556 16362 22568
rect 16960 22556 16988 22587
rect 17218 22584 17224 22636
rect 17276 22624 17282 22636
rect 17696 22624 17816 22628
rect 17276 22600 17816 22624
rect 17276 22596 17724 22600
rect 17276 22584 17282 22596
rect 17788 22565 17816 22600
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18472 22596 18521 22624
rect 18472 22584 18478 22596
rect 18509 22593 18521 22596
rect 18555 22624 18567 22627
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 18555 22596 19349 22624
rect 18555 22593 18567 22596
rect 18509 22587 18567 22593
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 20530 22584 20536 22636
rect 20588 22584 20594 22636
rect 21818 22584 21824 22636
rect 21876 22584 21882 22636
rect 24486 22584 24492 22636
rect 24544 22584 24550 22636
rect 16356 22528 16988 22556
rect 17681 22559 17739 22565
rect 16356 22516 16362 22528
rect 17681 22525 17693 22559
rect 17727 22525 17739 22559
rect 17681 22519 17739 22525
rect 17773 22559 17831 22565
rect 17773 22525 17785 22559
rect 17819 22525 17831 22559
rect 17773 22519 17831 22525
rect 15838 22448 15844 22500
rect 15896 22488 15902 22500
rect 16574 22488 16580 22500
rect 15896 22460 16580 22488
rect 15896 22448 15902 22460
rect 16574 22448 16580 22460
rect 16632 22448 16638 22500
rect 16850 22448 16856 22500
rect 16908 22488 16914 22500
rect 17586 22488 17592 22500
rect 16908 22460 17592 22488
rect 16908 22448 16914 22460
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 17696 22488 17724 22519
rect 19426 22516 19432 22568
rect 19484 22516 19490 22568
rect 19518 22516 19524 22568
rect 19576 22556 19582 22568
rect 19613 22559 19671 22565
rect 19613 22556 19625 22559
rect 19576 22528 19625 22556
rect 19576 22516 19582 22528
rect 19613 22525 19625 22528
rect 19659 22525 19671 22559
rect 20625 22559 20683 22565
rect 20625 22556 20637 22559
rect 19613 22519 19671 22525
rect 19727 22528 20637 22556
rect 17862 22488 17868 22500
rect 17696 22460 17868 22488
rect 17862 22448 17868 22460
rect 17920 22448 17926 22500
rect 18322 22448 18328 22500
rect 18380 22488 18386 22500
rect 19727 22488 19755 22528
rect 20625 22525 20637 22528
rect 20671 22525 20683 22559
rect 20625 22519 20683 22525
rect 20717 22559 20775 22565
rect 20717 22525 20729 22559
rect 20763 22525 20775 22559
rect 20717 22519 20775 22525
rect 20824 22528 22416 22556
rect 18380 22460 19755 22488
rect 18380 22448 18386 22460
rect 19794 22448 19800 22500
rect 19852 22488 19858 22500
rect 19978 22488 19984 22500
rect 19852 22460 19984 22488
rect 19852 22448 19858 22460
rect 19978 22448 19984 22460
rect 20036 22488 20042 22500
rect 20732 22488 20760 22519
rect 20036 22460 20760 22488
rect 20036 22448 20042 22460
rect 16390 22420 16396 22432
rect 13372 22392 16396 22420
rect 12897 22383 12955 22389
rect 16390 22380 16396 22392
rect 16448 22380 16454 22432
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 19518 22420 19524 22432
rect 17000 22392 19524 22420
rect 17000 22380 17006 22392
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20824 22420 20852 22528
rect 21637 22491 21695 22497
rect 21637 22457 21649 22491
rect 21683 22488 21695 22491
rect 22278 22488 22284 22500
rect 21683 22460 22284 22488
rect 21683 22457 21695 22460
rect 21637 22451 21695 22457
rect 22278 22448 22284 22460
rect 22336 22448 22342 22500
rect 22388 22488 22416 22528
rect 22462 22516 22468 22568
rect 22520 22516 22526 22568
rect 22649 22559 22707 22565
rect 22649 22525 22661 22559
rect 22695 22556 22707 22559
rect 22830 22556 22836 22568
rect 22695 22528 22836 22556
rect 22695 22525 22707 22528
rect 22649 22519 22707 22525
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 24581 22559 24639 22565
rect 24581 22556 24593 22559
rect 23676 22528 24593 22556
rect 22554 22488 22560 22500
rect 22388 22460 22560 22488
rect 22554 22448 22560 22460
rect 22612 22448 22618 22500
rect 23676 22432 23704 22528
rect 24581 22525 24593 22528
rect 24627 22525 24639 22559
rect 24581 22519 24639 22525
rect 24670 22516 24676 22568
rect 24728 22516 24734 22568
rect 20128 22392 20852 22420
rect 20128 22380 20134 22392
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21726 22420 21732 22432
rect 21048 22392 21732 22420
rect 21048 22380 21054 22392
rect 21726 22380 21732 22392
rect 21784 22380 21790 22432
rect 22002 22380 22008 22432
rect 22060 22380 22066 22432
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 23106 22420 23112 22432
rect 22244 22392 23112 22420
rect 22244 22380 22250 22392
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 23658 22380 23664 22432
rect 23716 22380 23722 22432
rect 24121 22423 24179 22429
rect 24121 22389 24133 22423
rect 24167 22420 24179 22423
rect 25038 22420 25044 22432
rect 24167 22392 25044 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 25038 22380 25044 22392
rect 25096 22380 25102 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 9953 22219 10011 22225
rect 9953 22216 9965 22219
rect 9824 22188 9965 22216
rect 9824 22176 9830 22188
rect 9953 22185 9965 22188
rect 9999 22185 10011 22219
rect 9953 22179 10011 22185
rect 10860 22219 10918 22225
rect 10860 22185 10872 22219
rect 10906 22216 10918 22219
rect 13630 22216 13636 22228
rect 10906 22188 13636 22216
rect 10906 22185 10918 22188
rect 10860 22179 10918 22185
rect 13630 22176 13636 22188
rect 13688 22216 13694 22228
rect 18598 22216 18604 22228
rect 13688 22188 16620 22216
rect 13688 22176 13694 22188
rect 2038 22108 2044 22160
rect 2096 22148 2102 22160
rect 2958 22148 2964 22160
rect 2096 22120 2964 22148
rect 2096 22108 2102 22120
rect 2958 22108 2964 22120
rect 3016 22108 3022 22160
rect 3602 22108 3608 22160
rect 3660 22148 3666 22160
rect 10502 22148 10508 22160
rect 3660 22120 10508 22148
rect 3660 22108 3666 22120
rect 10502 22108 10508 22120
rect 10560 22108 10566 22160
rect 11882 22108 11888 22160
rect 11940 22148 11946 22160
rect 11940 22120 12848 22148
rect 11940 22108 11946 22120
rect 2866 22040 2872 22092
rect 2924 22040 2930 22092
rect 6086 22040 6092 22092
rect 6144 22040 6150 22092
rect 8294 22040 8300 22092
rect 8352 22040 8358 22092
rect 9122 22040 9128 22092
rect 9180 22080 9186 22092
rect 9180 22052 10272 22080
rect 9180 22040 9186 22052
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 2271 21984 2774 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 2746 21876 2774 21984
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 4065 22015 4123 22021
rect 4065 22012 4077 22015
rect 3476 21984 4077 22012
rect 3476 21972 3482 21984
rect 4065 21981 4077 21984
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 4522 21972 4528 22024
rect 4580 22012 4586 22024
rect 4798 22012 4804 22024
rect 4580 21984 4804 22012
rect 4580 21972 4586 21984
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 4893 22015 4951 22021
rect 4893 21981 4905 22015
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 4249 21947 4307 21953
rect 4249 21913 4261 21947
rect 4295 21944 4307 21947
rect 4908 21944 4936 21975
rect 5534 21972 5540 22024
rect 5592 21972 5598 22024
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7466 22012 7472 22024
rect 7423 21984 7472 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 22012 9551 22015
rect 9539 21984 10088 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 9858 21944 9864 21956
rect 4295 21916 4844 21944
rect 4908 21916 9864 21944
rect 4295 21913 4307 21916
rect 4249 21907 4307 21913
rect 4522 21876 4528 21888
rect 2746 21848 4528 21876
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 4816 21876 4844 21916
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 7834 21876 7840 21888
rect 4816 21848 7840 21876
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 9309 21879 9367 21885
rect 9309 21876 9321 21879
rect 8904 21848 9321 21876
rect 8904 21836 8910 21848
rect 9309 21845 9321 21848
rect 9355 21845 9367 21879
rect 10060 21876 10088 21984
rect 10134 21972 10140 22024
rect 10192 21972 10198 22024
rect 10244 22012 10272 22052
rect 12158 22040 12164 22092
rect 12216 22080 12222 22092
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 12216 22052 12357 22080
rect 12216 22040 12222 22052
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12820 22080 12848 22120
rect 13262 22108 13268 22160
rect 13320 22148 13326 22160
rect 13722 22148 13728 22160
rect 13320 22120 13728 22148
rect 13320 22108 13326 22120
rect 13722 22108 13728 22120
rect 13780 22108 13786 22160
rect 13998 22108 14004 22160
rect 14056 22148 14062 22160
rect 14366 22148 14372 22160
rect 14056 22120 14372 22148
rect 14056 22108 14062 22120
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 14734 22108 14740 22160
rect 14792 22148 14798 22160
rect 14829 22151 14887 22157
rect 14829 22148 14841 22151
rect 14792 22120 14841 22148
rect 14792 22108 14798 22120
rect 14829 22117 14841 22120
rect 14875 22117 14887 22151
rect 14829 22111 14887 22117
rect 15194 22080 15200 22092
rect 12820 22052 15200 22080
rect 12345 22043 12403 22049
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15470 22040 15476 22092
rect 15528 22080 15534 22092
rect 16592 22089 16620 22188
rect 16684 22188 18604 22216
rect 16577 22083 16635 22089
rect 15528 22052 15700 22080
rect 15528 22040 15534 22052
rect 10594 22012 10600 22024
rect 10244 21984 10600 22012
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 12492 21984 13553 22012
rect 12492 21972 12498 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 15010 22012 15016 22024
rect 13780 21984 15016 22012
rect 13780 21972 13786 21984
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 15102 21972 15108 22024
rect 15160 22012 15166 22024
rect 15160 21984 15608 22012
rect 15160 21972 15166 21984
rect 11330 21904 11336 21956
rect 11388 21904 11394 21956
rect 14090 21944 14096 21956
rect 13372 21916 14096 21944
rect 13372 21876 13400 21916
rect 14090 21904 14096 21916
rect 14148 21904 14154 21956
rect 14642 21904 14648 21956
rect 14700 21904 14706 21956
rect 15378 21904 15384 21956
rect 15436 21904 15442 21956
rect 10060 21848 13400 21876
rect 9309 21839 9367 21845
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 13504 21848 15485 21876
rect 13504 21836 13510 21848
rect 15473 21845 15485 21848
rect 15519 21845 15531 21879
rect 15580 21876 15608 21984
rect 15672 21944 15700 22052
rect 16577 22049 16589 22083
rect 16623 22049 16635 22083
rect 16577 22043 16635 22049
rect 16390 21972 16396 22024
rect 16448 22012 16454 22024
rect 16684 22012 16712 22188
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 18874 22176 18880 22228
rect 18932 22216 18938 22228
rect 20806 22216 20812 22228
rect 18932 22188 20812 22216
rect 18932 22176 18938 22188
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 21726 22176 21732 22228
rect 21784 22216 21790 22228
rect 21910 22216 21916 22228
rect 21784 22188 21916 22216
rect 21784 22176 21790 22188
rect 21910 22176 21916 22188
rect 21968 22176 21974 22228
rect 17313 22151 17371 22157
rect 17313 22117 17325 22151
rect 17359 22117 17371 22151
rect 17313 22111 17371 22117
rect 17880 22120 18644 22148
rect 16448 21984 16712 22012
rect 16448 21972 16454 21984
rect 17328 21944 17356 22111
rect 17402 22040 17408 22092
rect 17460 22080 17466 22092
rect 17880 22080 17908 22120
rect 17460 22052 17908 22080
rect 17957 22083 18015 22089
rect 17460 22040 17466 22052
rect 17957 22049 17969 22083
rect 18003 22080 18015 22083
rect 18506 22080 18512 22092
rect 18003 22052 18512 22080
rect 18003 22049 18015 22052
rect 17957 22043 18015 22049
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 18616 22080 18644 22120
rect 22278 22108 22284 22160
rect 22336 22148 22342 22160
rect 23290 22148 23296 22160
rect 22336 22120 23296 22148
rect 22336 22108 22342 22120
rect 18616 22052 19840 22080
rect 19812 22021 19840 22052
rect 20070 22040 20076 22092
rect 20128 22040 20134 22092
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 22094 22080 22100 22092
rect 20487 22052 22100 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 22094 22040 22100 22052
rect 22152 22040 22158 22092
rect 22189 22083 22247 22089
rect 22189 22049 22201 22083
rect 22235 22080 22247 22083
rect 22370 22080 22376 22092
rect 22235 22052 22376 22080
rect 22235 22049 22247 22052
rect 22189 22043 22247 22049
rect 22370 22040 22376 22052
rect 22428 22040 22434 22092
rect 22480 22089 22508 22120
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 23474 22108 23480 22160
rect 23532 22148 23538 22160
rect 24486 22148 24492 22160
rect 23532 22120 24492 22148
rect 23532 22108 23538 22120
rect 24486 22108 24492 22120
rect 24544 22108 24550 22160
rect 25130 22108 25136 22160
rect 25188 22148 25194 22160
rect 25188 22120 25268 22148
rect 25188 22108 25194 22120
rect 25240 22089 25268 22120
rect 22465 22083 22523 22089
rect 22465 22049 22477 22083
rect 22511 22049 22523 22083
rect 22465 22043 22523 22049
rect 25225 22083 25283 22089
rect 25225 22049 25237 22083
rect 25271 22080 25283 22083
rect 25271 22052 25305 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 25406 22040 25412 22092
rect 25464 22040 25470 22092
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 22012 17831 22015
rect 19797 22015 19855 22021
rect 17819 21984 19472 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 17862 21944 17868 21956
rect 15672 21916 17356 21944
rect 17420 21916 17868 21944
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 15580 21848 16037 21876
rect 15473 21839 15531 21845
rect 16025 21845 16037 21848
rect 16071 21845 16083 21879
rect 16025 21839 16083 21845
rect 16114 21836 16120 21888
rect 16172 21876 16178 21888
rect 16393 21879 16451 21885
rect 16393 21876 16405 21879
rect 16172 21848 16405 21876
rect 16172 21836 16178 21848
rect 16393 21845 16405 21848
rect 16439 21845 16451 21879
rect 16393 21839 16451 21845
rect 16485 21879 16543 21885
rect 16485 21845 16497 21879
rect 16531 21876 16543 21879
rect 16758 21876 16764 21888
rect 16531 21848 16764 21876
rect 16531 21845 16543 21848
rect 16485 21839 16543 21845
rect 16758 21836 16764 21848
rect 16816 21876 16822 21888
rect 17420 21876 17448 21916
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 18598 21904 18604 21956
rect 18656 21904 18662 21956
rect 16816 21848 17448 21876
rect 16816 21836 16822 21848
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 18690 21836 18696 21888
rect 18748 21836 18754 21888
rect 19444 21885 19472 21984
rect 19797 21981 19809 22015
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 22741 22015 22799 22021
rect 22741 21981 22753 22015
rect 22787 22012 22799 22015
rect 23290 22012 23296 22024
rect 22787 21984 23296 22012
rect 22787 21981 22799 21984
rect 22741 21975 22799 21981
rect 23290 21972 23296 21984
rect 23348 22012 23354 22024
rect 25424 22012 25452 22040
rect 23348 21984 25452 22012
rect 23348 21972 23354 21984
rect 20717 21947 20775 21953
rect 20717 21913 20729 21947
rect 20763 21944 20775 21947
rect 20990 21944 20996 21956
rect 20763 21916 20996 21944
rect 20763 21913 20775 21916
rect 20717 21907 20775 21913
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 21726 21904 21732 21956
rect 21784 21904 21790 21956
rect 25041 21947 25099 21953
rect 25041 21944 25053 21947
rect 23768 21916 25053 21944
rect 19429 21879 19487 21885
rect 19429 21845 19441 21879
rect 19475 21845 19487 21879
rect 19429 21839 19487 21845
rect 19702 21836 19708 21888
rect 19760 21876 19766 21888
rect 19889 21879 19947 21885
rect 19889 21876 19901 21879
rect 19760 21848 19901 21876
rect 19760 21836 19766 21848
rect 19889 21845 19901 21848
rect 19935 21845 19947 21879
rect 19889 21839 19947 21845
rect 21358 21836 21364 21888
rect 21416 21876 21422 21888
rect 23474 21876 23480 21888
rect 21416 21848 23480 21876
rect 21416 21836 21422 21848
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 23768 21885 23796 21916
rect 25041 21913 25053 21916
rect 25087 21913 25099 21947
rect 25041 21907 25099 21913
rect 23753 21879 23811 21885
rect 23753 21876 23765 21879
rect 23624 21848 23765 21876
rect 23624 21836 23630 21848
rect 23753 21845 23765 21848
rect 23799 21845 23811 21879
rect 23753 21839 23811 21845
rect 24578 21836 24584 21888
rect 24636 21836 24642 21888
rect 24949 21879 25007 21885
rect 24949 21845 24961 21879
rect 24995 21876 25007 21879
rect 25314 21876 25320 21888
rect 24995 21848 25320 21876
rect 24995 21845 25007 21848
rect 24949 21839 25007 21845
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 2774 21672 2780 21684
rect 2746 21632 2780 21672
rect 2832 21632 2838 21684
rect 2884 21644 12020 21672
rect 1673 21607 1731 21613
rect 1673 21573 1685 21607
rect 1719 21604 1731 21607
rect 2746 21604 2774 21632
rect 1719 21576 2774 21604
rect 1719 21573 1731 21576
rect 1673 21567 1731 21573
rect 1857 21471 1915 21477
rect 1857 21437 1869 21471
rect 1903 21468 1915 21471
rect 2884 21468 2912 21644
rect 6730 21604 6736 21616
rect 2976 21576 6736 21604
rect 2976 21545 3004 21576
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 10870 21604 10876 21616
rect 10626 21576 10876 21604
rect 10870 21564 10876 21576
rect 10928 21604 10934 21616
rect 11330 21604 11336 21616
rect 10928 21576 11336 21604
rect 10928 21564 10934 21576
rect 11330 21564 11336 21576
rect 11388 21564 11394 21616
rect 11992 21604 12020 21644
rect 12066 21632 12072 21684
rect 12124 21632 12130 21684
rect 12434 21632 12440 21684
rect 12492 21632 12498 21684
rect 14550 21672 14556 21684
rect 13563 21644 14556 21672
rect 13262 21604 13268 21616
rect 11992 21576 13268 21604
rect 13262 21564 13268 21576
rect 13320 21564 13326 21616
rect 13563 21613 13591 21644
rect 14550 21632 14556 21644
rect 14608 21632 14614 21684
rect 15473 21675 15531 21681
rect 15473 21641 15485 21675
rect 15519 21672 15531 21675
rect 16022 21672 16028 21684
rect 15519 21644 16028 21672
rect 15519 21641 15531 21644
rect 15473 21635 15531 21641
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 17034 21632 17040 21684
rect 17092 21672 17098 21684
rect 17402 21672 17408 21684
rect 17092 21644 17408 21672
rect 17092 21632 17098 21644
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 17678 21632 17684 21684
rect 17736 21672 17742 21684
rect 17736 21644 19932 21672
rect 17736 21632 17742 21644
rect 13541 21607 13599 21613
rect 13541 21573 13553 21607
rect 13587 21573 13599 21607
rect 13541 21567 13599 21573
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 17497 21607 17555 21613
rect 17497 21604 17509 21607
rect 13872 21576 14030 21604
rect 14844 21576 17509 21604
rect 13872 21564 13878 21576
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 8570 21536 8576 21548
rect 7515 21508 8576 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 8570 21496 8576 21508
rect 8628 21496 8634 21548
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12216 21508 12664 21536
rect 12216 21496 12222 21508
rect 1903 21440 2912 21468
rect 1903 21437 1915 21440
rect 1857 21431 1915 21437
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 4982 21428 4988 21480
rect 5040 21468 5046 21480
rect 5077 21471 5135 21477
rect 5077 21468 5089 21471
rect 5040 21440 5089 21468
rect 5040 21428 5046 21440
rect 5077 21437 5089 21440
rect 5123 21437 5135 21471
rect 5077 21431 5135 21437
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 7745 21471 7803 21477
rect 7745 21468 7757 21471
rect 7248 21440 7757 21468
rect 7248 21428 7254 21440
rect 7745 21437 7757 21440
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 9122 21428 9128 21480
rect 9180 21428 9186 21480
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 11146 21468 11152 21480
rect 9447 21440 11152 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 12526 21428 12532 21480
rect 12584 21428 12590 21480
rect 12636 21477 12664 21508
rect 12621 21471 12679 21477
rect 12621 21437 12633 21471
rect 12667 21437 12679 21471
rect 12621 21431 12679 21437
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 13265 21471 13323 21477
rect 13265 21468 13277 21471
rect 12768 21440 13277 21468
rect 12768 21428 12774 21440
rect 13265 21437 13277 21440
rect 13311 21437 13323 21471
rect 14844 21468 14872 21576
rect 17497 21573 17509 21576
rect 17543 21573 17555 21607
rect 18782 21604 18788 21616
rect 17497 21567 17555 21573
rect 18248 21576 18788 21604
rect 15010 21496 15016 21548
rect 15068 21536 15074 21548
rect 15286 21536 15292 21548
rect 15068 21508 15292 21536
rect 15068 21496 15074 21508
rect 15286 21496 15292 21508
rect 15344 21536 15350 21548
rect 15841 21539 15899 21545
rect 15841 21536 15853 21539
rect 15344 21508 15853 21536
rect 15344 21496 15350 21508
rect 15841 21505 15853 21508
rect 15887 21505 15899 21539
rect 15841 21499 15899 21505
rect 17402 21496 17408 21548
rect 17460 21496 17466 21548
rect 17770 21496 17776 21548
rect 17828 21536 17834 21548
rect 18248 21545 18276 21576
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 19904 21604 19932 21644
rect 19978 21632 19984 21684
rect 20036 21632 20042 21684
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 23566 21672 23572 21684
rect 20312 21644 23572 21672
rect 20312 21632 20318 21644
rect 23566 21632 23572 21644
rect 23624 21632 23630 21684
rect 24026 21632 24032 21684
rect 24084 21632 24090 21684
rect 25038 21632 25044 21684
rect 25096 21632 25102 21684
rect 22646 21604 22652 21616
rect 19904 21576 22652 21604
rect 22646 21564 22652 21576
rect 22704 21564 22710 21616
rect 23842 21604 23848 21616
rect 23782 21576 23848 21604
rect 23842 21564 23848 21576
rect 23900 21564 23906 21616
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 17828 21508 18245 21536
rect 17828 21496 17834 21508
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 19610 21496 19616 21548
rect 19668 21496 19674 21548
rect 20806 21496 20812 21548
rect 20864 21536 20870 21548
rect 21358 21536 21364 21548
rect 20864 21508 21364 21536
rect 20864 21496 20870 21508
rect 21358 21496 21364 21508
rect 21416 21496 21422 21548
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21536 25007 21539
rect 25038 21536 25044 21548
rect 24995 21508 25044 21536
rect 24995 21505 25007 21508
rect 24949 21499 25007 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 13265 21431 13323 21437
rect 13372 21440 14872 21468
rect 10410 21360 10416 21412
rect 10468 21400 10474 21412
rect 13372 21400 13400 21440
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 15528 21440 15945 21468
rect 15528 21428 15534 21440
rect 15933 21437 15945 21440
rect 15979 21468 15991 21471
rect 16022 21468 16028 21480
rect 15979 21440 16028 21468
rect 15979 21437 15991 21440
rect 15933 21431 15991 21437
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 16117 21471 16175 21477
rect 16117 21437 16129 21471
rect 16163 21468 16175 21471
rect 17494 21468 17500 21480
rect 16163 21440 17500 21468
rect 16163 21437 16175 21440
rect 16117 21431 16175 21437
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 17678 21428 17684 21480
rect 17736 21428 17742 21480
rect 18506 21428 18512 21480
rect 18564 21428 18570 21480
rect 18874 21428 18880 21480
rect 18932 21468 18938 21480
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 18932 21440 20913 21468
rect 18932 21428 18938 21440
rect 20901 21437 20913 21440
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 21085 21471 21143 21477
rect 21085 21437 21097 21471
rect 21131 21468 21143 21471
rect 21266 21468 21272 21480
rect 21131 21440 21272 21468
rect 21131 21437 21143 21440
rect 21085 21431 21143 21437
rect 21266 21428 21272 21440
rect 21324 21428 21330 21480
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22281 21471 22339 21477
rect 22281 21468 22293 21471
rect 22152 21440 22293 21468
rect 22152 21428 22158 21440
rect 22281 21437 22293 21440
rect 22327 21437 22339 21471
rect 22554 21468 22560 21480
rect 22281 21431 22339 21437
rect 22388 21440 22560 21468
rect 10468 21372 13400 21400
rect 14568 21372 15148 21400
rect 10468 21360 10474 21372
rect 6825 21335 6883 21341
rect 6825 21301 6837 21335
rect 6871 21332 6883 21335
rect 10134 21332 10140 21344
rect 6871 21304 10140 21332
rect 6871 21301 6883 21304
rect 6825 21295 6883 21301
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 10873 21335 10931 21341
rect 10873 21332 10885 21335
rect 10744 21304 10885 21332
rect 10744 21292 10750 21304
rect 10873 21301 10885 21304
rect 10919 21301 10931 21335
rect 10873 21295 10931 21301
rect 10962 21292 10968 21344
rect 11020 21332 11026 21344
rect 12434 21332 12440 21344
rect 11020 21304 12440 21332
rect 11020 21292 11026 21304
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 12526 21292 12532 21344
rect 12584 21332 12590 21344
rect 13722 21332 13728 21344
rect 12584 21304 13728 21332
rect 12584 21292 12590 21304
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 14568 21332 14596 21372
rect 14148 21304 14596 21332
rect 14148 21292 14154 21304
rect 15010 21292 15016 21344
rect 15068 21292 15074 21344
rect 15120 21332 15148 21372
rect 15378 21360 15384 21412
rect 15436 21400 15442 21412
rect 18046 21400 18052 21412
rect 15436 21372 18052 21400
rect 15436 21360 15442 21372
rect 18046 21360 18052 21372
rect 18104 21360 18110 21412
rect 22388 21400 22416 21440
rect 22554 21428 22560 21440
rect 22612 21428 22618 21480
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 24305 21471 24363 21477
rect 24305 21468 24317 21471
rect 22704 21440 24317 21468
rect 22704 21428 22710 21440
rect 24305 21437 24317 21440
rect 24351 21437 24363 21471
rect 24305 21431 24363 21437
rect 25133 21471 25191 21477
rect 25133 21437 25145 21471
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 19536 21372 22416 21400
rect 16666 21332 16672 21344
rect 15120 21304 16672 21332
rect 16666 21292 16672 21304
rect 16724 21292 16730 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 19536 21332 19564 21372
rect 23750 21360 23756 21412
rect 23808 21400 23814 21412
rect 25148 21400 25176 21431
rect 23808 21372 25176 21400
rect 23808 21360 23814 21372
rect 17083 21304 19564 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 20438 21292 20444 21344
rect 20496 21292 20502 21344
rect 20990 21292 20996 21344
rect 21048 21332 21054 21344
rect 22002 21332 22008 21344
rect 21048 21304 22008 21332
rect 21048 21292 21054 21304
rect 22002 21292 22008 21304
rect 22060 21332 22066 21344
rect 22370 21332 22376 21344
rect 22060 21304 22376 21332
rect 22060 21292 22066 21304
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 22544 21335 22602 21341
rect 22544 21301 22556 21335
rect 22590 21332 22602 21335
rect 23658 21332 23664 21344
rect 22590 21304 23664 21332
rect 22590 21301 22602 21304
rect 22544 21295 22602 21301
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 24581 21335 24639 21341
rect 24581 21301 24593 21335
rect 24627 21332 24639 21335
rect 25682 21332 25688 21344
rect 24627 21304 25688 21332
rect 24627 21301 24639 21304
rect 24581 21295 24639 21301
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 2038 21088 2044 21140
rect 2096 21128 2102 21140
rect 7742 21128 7748 21140
rect 2096 21100 7748 21128
rect 2096 21088 2102 21100
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 12897 21131 12955 21137
rect 10520 21100 12848 21128
rect 2774 21020 2780 21072
rect 2832 21060 2838 21072
rect 2832 21032 2912 21060
rect 2832 21020 2838 21032
rect 2884 21001 2912 21032
rect 6914 21020 6920 21072
rect 6972 21020 6978 21072
rect 7006 21020 7012 21072
rect 7064 21060 7070 21072
rect 7064 21032 7512 21060
rect 7064 21020 7070 21032
rect 2869 20995 2927 21001
rect 2240 20964 2774 20992
rect 2240 20933 2268 20964
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 2746 20856 2774 20964
rect 2869 20961 2881 20995
rect 2915 20961 2927 20995
rect 2869 20955 2927 20961
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 6932 20992 6960 21020
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 6932 20964 7389 20992
rect 4433 20955 4491 20961
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 7484 20992 7512 21032
rect 10413 20995 10471 21001
rect 7484 20964 10364 20992
rect 7377 20955 7435 20961
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 5718 20924 5724 20936
rect 4111 20896 5724 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20924 6055 20927
rect 6546 20924 6552 20936
rect 6043 20896 6552 20924
rect 6043 20893 6055 20896
rect 5997 20887 6055 20893
rect 6546 20884 6552 20896
rect 6604 20884 6610 20936
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7650 20924 7656 20936
rect 7147 20896 7656 20924
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 10336 20924 10364 20964
rect 10413 20961 10425 20995
rect 10459 20992 10471 20995
rect 10520 20992 10548 21100
rect 12434 21020 12440 21072
rect 12492 21060 12498 21072
rect 12820 21060 12848 21100
rect 12897 21097 12909 21131
rect 12943 21128 12955 21131
rect 13630 21128 13636 21140
rect 12943 21100 13636 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 15473 21131 15531 21137
rect 15473 21128 15485 21131
rect 13924 21100 15485 21128
rect 13924 21060 13952 21100
rect 15473 21097 15485 21100
rect 15519 21097 15531 21131
rect 15473 21091 15531 21097
rect 16850 21088 16856 21140
rect 16908 21088 16914 21140
rect 16942 21088 16948 21140
rect 17000 21128 17006 21140
rect 19613 21131 19671 21137
rect 17000 21100 19012 21128
rect 17000 21088 17006 21100
rect 12492 21032 12756 21060
rect 12820 21032 13952 21060
rect 12492 21020 12498 21032
rect 10459 20964 10548 20992
rect 10597 20995 10655 21001
rect 10459 20961 10471 20964
rect 10413 20955 10471 20961
rect 10597 20961 10609 20995
rect 10643 20992 10655 20995
rect 10686 20992 10692 21004
rect 10643 20964 10692 20992
rect 10643 20961 10655 20964
rect 10597 20955 10655 20961
rect 10686 20952 10692 20964
rect 10744 20952 10750 21004
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20992 11207 20995
rect 12728 20992 12756 21032
rect 14274 21020 14280 21072
rect 14332 21020 14338 21072
rect 17497 21063 17555 21069
rect 17497 21060 17509 21063
rect 14752 21032 17509 21060
rect 14090 20992 14096 21004
rect 11195 20964 12664 20992
rect 12728 20964 14096 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 10962 20924 10968 20936
rect 10336 20896 10968 20924
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 6454 20856 6460 20868
rect 2746 20828 6460 20856
rect 6454 20816 6460 20828
rect 6512 20816 6518 20868
rect 10410 20856 10416 20868
rect 9140 20828 10416 20856
rect 5810 20748 5816 20800
rect 5868 20748 5874 20800
rect 9140 20797 9168 20828
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 10594 20816 10600 20868
rect 10652 20856 10658 20868
rect 11164 20856 11192 20955
rect 12636 20924 12664 20964
rect 14090 20952 14096 20964
rect 14148 20952 14154 21004
rect 14752 21001 14780 21032
rect 17497 21029 17509 21032
rect 17543 21029 17555 21063
rect 18874 21060 18880 21072
rect 17497 21023 17555 21029
rect 18156 21032 18880 21060
rect 14737 20995 14795 21001
rect 14737 20961 14749 20995
rect 14783 20961 14795 20995
rect 14737 20955 14795 20961
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 15102 20992 15108 21004
rect 14967 20964 15108 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 15102 20952 15108 20964
rect 15160 20952 15166 21004
rect 15194 20952 15200 21004
rect 15252 20992 15258 21004
rect 16025 20995 16083 21001
rect 16025 20992 16037 20995
rect 15252 20964 16037 20992
rect 15252 20952 15258 20964
rect 16025 20961 16037 20964
rect 16071 20961 16083 20995
rect 18049 20995 18107 21001
rect 18049 20992 18061 20995
rect 16025 20955 16083 20961
rect 16132 20964 18061 20992
rect 12710 20924 12716 20936
rect 12636 20896 12716 20924
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 12802 20884 12808 20936
rect 12860 20924 12866 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 12860 20896 13553 20924
rect 12860 20884 12866 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 14645 20927 14703 20933
rect 14645 20924 14657 20927
rect 14516 20896 14657 20924
rect 14516 20884 14522 20896
rect 14645 20893 14657 20896
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 15010 20884 15016 20936
rect 15068 20924 15074 20936
rect 16132 20924 16160 20964
rect 18049 20961 18061 20964
rect 18095 20961 18107 20995
rect 18049 20955 18107 20961
rect 18156 20924 18184 21032
rect 18874 21020 18880 21032
rect 18932 21020 18938 21072
rect 18984 21060 19012 21100
rect 19613 21097 19625 21131
rect 19659 21128 19671 21131
rect 20806 21128 20812 21140
rect 19659 21100 20812 21128
rect 19659 21097 19671 21100
rect 19613 21091 19671 21097
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 22370 21088 22376 21140
rect 22428 21128 22434 21140
rect 23750 21128 23756 21140
rect 22428 21100 23756 21128
rect 22428 21088 22434 21100
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 24210 21088 24216 21140
rect 24268 21088 24274 21140
rect 20254 21060 20260 21072
rect 18984 21032 20260 21060
rect 20254 21020 20260 21032
rect 20312 21020 20318 21072
rect 21726 21020 21732 21072
rect 21784 21060 21790 21072
rect 21784 21032 21864 21060
rect 21784 21020 21790 21032
rect 18782 20952 18788 21004
rect 18840 20992 18846 21004
rect 20349 20995 20407 21001
rect 20349 20992 20361 20995
rect 18840 20964 20361 20992
rect 18840 20952 18846 20964
rect 20349 20961 20361 20964
rect 20395 20961 20407 20995
rect 20349 20955 20407 20961
rect 20625 20995 20683 21001
rect 20625 20961 20637 20995
rect 20671 20992 20683 20995
rect 20714 20992 20720 21004
rect 20671 20964 20720 20992
rect 20671 20961 20683 20964
rect 20625 20955 20683 20961
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 15068 20896 16160 20924
rect 16224 20896 18184 20924
rect 18877 20927 18935 20933
rect 15068 20884 15074 20896
rect 10652 20828 11192 20856
rect 11425 20859 11483 20865
rect 10652 20816 10658 20828
rect 11425 20825 11437 20859
rect 11471 20825 11483 20859
rect 13630 20856 13636 20868
rect 12650 20828 13636 20856
rect 11425 20819 11483 20825
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20757 9183 20791
rect 9125 20751 9183 20757
rect 9950 20748 9956 20800
rect 10008 20748 10014 20800
rect 10134 20748 10140 20800
rect 10192 20788 10198 20800
rect 10321 20791 10379 20797
rect 10321 20788 10333 20791
rect 10192 20760 10333 20788
rect 10192 20748 10198 20760
rect 10321 20757 10333 20760
rect 10367 20757 10379 20791
rect 11440 20788 11468 20819
rect 13630 20816 13636 20828
rect 13688 20856 13694 20868
rect 13814 20856 13820 20868
rect 13688 20828 13820 20856
rect 13688 20816 13694 20828
rect 13814 20816 13820 20828
rect 13872 20856 13878 20868
rect 14274 20856 14280 20868
rect 13872 20828 14280 20856
rect 13872 20816 13878 20828
rect 14274 20816 14280 20828
rect 14332 20816 14338 20868
rect 15470 20816 15476 20868
rect 15528 20856 15534 20868
rect 16224 20856 16252 20896
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 19794 20924 19800 20936
rect 18923 20896 19800 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 21836 20924 21864 21032
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 22097 21063 22155 21069
rect 22097 21060 22109 21063
rect 22060 21032 22109 21060
rect 22060 21020 22066 21032
rect 22097 21029 22109 21032
rect 22143 21029 22155 21063
rect 22097 21023 22155 21029
rect 21910 20952 21916 21004
rect 21968 20992 21974 21004
rect 22186 20992 22192 21004
rect 21968 20964 22192 20992
rect 21968 20952 21974 20964
rect 22186 20952 22192 20964
rect 22244 20952 22250 21004
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 23382 20992 23388 21004
rect 22787 20964 23388 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 23474 20952 23480 21004
rect 23532 20992 23538 21004
rect 24949 20995 25007 21001
rect 24949 20992 24961 20995
rect 23532 20964 24961 20992
rect 23532 20952 23538 20964
rect 24949 20961 24961 20964
rect 24995 20961 25007 20995
rect 24949 20955 25007 20961
rect 21836 20896 21956 20924
rect 15528 20828 16252 20856
rect 15528 20816 15534 20828
rect 16758 20816 16764 20868
rect 16816 20816 16822 20868
rect 17126 20856 17132 20868
rect 16868 20828 17132 20856
rect 12158 20788 12164 20800
rect 11440 20760 12164 20788
rect 10321 20751 10379 20757
rect 12158 20748 12164 20760
rect 12216 20788 12222 20800
rect 13354 20788 13360 20800
rect 12216 20760 13360 20788
rect 12216 20748 12222 20760
rect 13354 20748 13360 20760
rect 13412 20748 13418 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 15841 20791 15899 20797
rect 15841 20788 15853 20791
rect 14792 20760 15853 20788
rect 14792 20748 14798 20760
rect 15841 20757 15853 20760
rect 15887 20757 15899 20791
rect 15841 20751 15899 20757
rect 15933 20791 15991 20797
rect 15933 20757 15945 20791
rect 15979 20788 15991 20791
rect 16666 20788 16672 20800
rect 15979 20760 16672 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16666 20748 16672 20760
rect 16724 20788 16730 20800
rect 16868 20788 16896 20828
rect 17126 20816 17132 20828
rect 17184 20856 17190 20868
rect 17957 20859 18015 20865
rect 17957 20856 17969 20859
rect 17184 20828 17969 20856
rect 17184 20816 17190 20828
rect 17957 20825 17969 20828
rect 18003 20856 18015 20859
rect 18322 20856 18328 20868
rect 18003 20828 18328 20856
rect 18003 20825 18015 20828
rect 17957 20819 18015 20825
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 19610 20856 19616 20868
rect 19392 20828 19616 20856
rect 19392 20816 19398 20828
rect 19610 20816 19616 20828
rect 19668 20856 19674 20868
rect 21082 20856 21088 20868
rect 19668 20828 21088 20856
rect 19668 20816 19674 20828
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 21928 20856 21956 20896
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22152 20896 22477 20924
rect 22152 20884 22158 20896
rect 22465 20893 22477 20896
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 23842 20884 23848 20936
rect 23900 20924 23906 20936
rect 24302 20924 24308 20936
rect 23900 20896 24308 20924
rect 23900 20884 23906 20896
rect 24302 20884 24308 20896
rect 24360 20884 24366 20936
rect 24486 20884 24492 20936
rect 24544 20924 24550 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24544 20896 24777 20924
rect 24544 20884 24550 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 22646 20856 22652 20868
rect 21850 20828 22652 20856
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 24026 20816 24032 20868
rect 24084 20856 24090 20868
rect 24857 20859 24915 20865
rect 24857 20856 24869 20859
rect 24084 20828 24869 20856
rect 24084 20816 24090 20828
rect 24857 20825 24869 20828
rect 24903 20825 24915 20859
rect 24857 20819 24915 20825
rect 16724 20760 16896 20788
rect 16724 20748 16730 20760
rect 16942 20748 16948 20800
rect 17000 20788 17006 20800
rect 17865 20791 17923 20797
rect 17865 20788 17877 20791
rect 17000 20760 17877 20788
rect 17000 20748 17006 20760
rect 17865 20757 17877 20760
rect 17911 20757 17923 20791
rect 17865 20751 17923 20757
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 18690 20788 18696 20800
rect 18104 20760 18696 20788
rect 18104 20748 18110 20760
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 20622 20748 20628 20800
rect 20680 20788 20686 20800
rect 23382 20788 23388 20800
rect 20680 20760 23388 20788
rect 20680 20748 20686 20760
rect 23382 20748 23388 20760
rect 23440 20748 23446 20800
rect 24394 20748 24400 20800
rect 24452 20748 24458 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 8386 20584 8392 20596
rect 1872 20556 8392 20584
rect 1872 20457 1900 20556
rect 8386 20544 8392 20556
rect 8444 20544 8450 20596
rect 8588 20556 10732 20584
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20417 1915 20451
rect 1857 20411 1915 20417
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 3007 20420 5948 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 1581 20383 1639 20389
rect 1581 20349 1593 20383
rect 1627 20349 1639 20383
rect 1581 20343 1639 20349
rect 1596 20312 1624 20343
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 5920 20380 5948 20420
rect 5994 20408 6000 20460
rect 6052 20408 6058 20460
rect 7098 20408 7104 20460
rect 7156 20408 7162 20460
rect 8588 20457 8616 20556
rect 9582 20516 9588 20528
rect 8864 20488 9588 20516
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 6914 20380 6920 20392
rect 5920 20352 6920 20380
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7377 20383 7435 20389
rect 7377 20349 7389 20383
rect 7423 20380 7435 20383
rect 8864 20380 8892 20488
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 10704 20516 10732 20556
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 12250 20584 12256 20596
rect 10836 20556 12256 20584
rect 10836 20544 10842 20556
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12802 20584 12808 20596
rect 12483 20556 12808 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12802 20544 12808 20556
rect 12860 20544 12866 20596
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 14826 20584 14832 20596
rect 13504 20556 14832 20584
rect 13504 20544 13510 20556
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15252 20556 15945 20584
rect 15252 20544 15258 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 18693 20587 18751 20593
rect 18693 20584 18705 20587
rect 18564 20556 18705 20584
rect 18564 20544 18570 20556
rect 18693 20553 18705 20556
rect 18739 20553 18751 20587
rect 18693 20547 18751 20553
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 22373 20587 22431 20593
rect 22373 20584 22385 20587
rect 20864 20556 22385 20584
rect 20864 20544 20870 20556
rect 22373 20553 22385 20556
rect 22419 20553 22431 20587
rect 22373 20547 22431 20553
rect 22465 20587 22523 20593
rect 22465 20553 22477 20587
rect 22511 20584 22523 20587
rect 23290 20584 23296 20596
rect 22511 20556 23296 20584
rect 22511 20553 22523 20556
rect 22465 20547 22523 20553
rect 11514 20516 11520 20528
rect 10704 20488 11520 20516
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 14274 20476 14280 20528
rect 14332 20476 14338 20528
rect 19610 20516 19616 20528
rect 18446 20488 19616 20516
rect 18524 20460 18552 20488
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 21082 20516 21088 20528
rect 20746 20488 21088 20516
rect 21082 20476 21088 20488
rect 21140 20476 21146 20528
rect 10594 20448 10600 20460
rect 10442 20420 10600 20448
rect 10594 20408 10600 20420
rect 10652 20448 10658 20460
rect 10870 20448 10876 20460
rect 10652 20420 10876 20448
rect 10652 20408 10658 20420
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 13446 20448 13452 20460
rect 11020 20420 13452 20448
rect 11020 20408 11026 20420
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 15930 20448 15936 20460
rect 15887 20420 15936 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 19242 20448 19248 20460
rect 18840 20420 19248 20448
rect 18840 20408 18846 20420
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 22480 20392 22508 20547
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 23198 20476 23204 20528
rect 23256 20476 23262 20528
rect 24302 20476 24308 20528
rect 24360 20476 24366 20528
rect 7423 20352 8892 20380
rect 7423 20349 7435 20352
rect 7377 20343 7435 20349
rect 9030 20340 9036 20392
rect 9088 20340 9094 20392
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 10686 20380 10692 20392
rect 9355 20352 10692 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 3694 20312 3700 20324
rect 1596 20284 3700 20312
rect 3694 20272 3700 20284
rect 3752 20272 3758 20324
rect 4709 20315 4767 20321
rect 4709 20281 4721 20315
rect 4755 20312 4767 20315
rect 5353 20315 5411 20321
rect 5353 20312 5365 20315
rect 4755 20284 5365 20312
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 5353 20281 5365 20284
rect 5399 20312 5411 20315
rect 8938 20312 8944 20324
rect 5399 20284 8944 20312
rect 5399 20281 5411 20284
rect 5353 20275 5411 20281
rect 8938 20272 8944 20284
rect 8996 20272 9002 20324
rect 12069 20315 12127 20321
rect 12069 20312 12081 20315
rect 10336 20284 12081 20312
rect 5813 20247 5871 20253
rect 5813 20213 5825 20247
rect 5859 20244 5871 20247
rect 7834 20244 7840 20256
rect 5859 20216 7840 20244
rect 5859 20213 5871 20216
rect 5813 20207 5871 20213
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 8386 20204 8392 20256
rect 8444 20204 8450 20256
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 10336 20244 10364 20284
rect 12069 20281 12081 20284
rect 12115 20281 12127 20315
rect 12069 20275 12127 20281
rect 8536 20216 10364 20244
rect 8536 20204 8542 20216
rect 10686 20204 10692 20256
rect 10744 20244 10750 20256
rect 10781 20247 10839 20253
rect 10781 20244 10793 20247
rect 10744 20216 10793 20244
rect 10744 20204 10750 20216
rect 10781 20213 10793 20216
rect 10827 20213 10839 20247
rect 12544 20244 12572 20343
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 15010 20380 15016 20392
rect 13863 20352 15016 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 16298 20380 16304 20392
rect 15252 20352 16304 20380
rect 15252 20340 15258 20352
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 16482 20340 16488 20392
rect 16540 20380 16546 20392
rect 16945 20383 17003 20389
rect 16945 20380 16957 20383
rect 16540 20352 16957 20380
rect 16540 20340 16546 20352
rect 16945 20349 16957 20352
rect 16991 20349 17003 20383
rect 16945 20343 17003 20349
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17276 20352 18276 20380
rect 17276 20340 17282 20352
rect 14918 20272 14924 20324
rect 14976 20312 14982 20324
rect 14976 20284 15424 20312
rect 14976 20272 14982 20284
rect 15010 20244 15016 20256
rect 12544 20216 15016 20244
rect 10781 20207 10839 20213
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 15160 20216 15301 20244
rect 15160 20204 15166 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15396 20244 15424 20284
rect 17954 20244 17960 20256
rect 15396 20216 17960 20244
rect 15289 20207 15347 20213
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 18248 20244 18276 20352
rect 19518 20340 19524 20392
rect 19576 20340 19582 20392
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20772 20352 21005 20380
rect 20772 20340 20778 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 22462 20380 22468 20392
rect 20993 20343 21051 20349
rect 21100 20352 22468 20380
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 21100 20312 21128 20352
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 22572 20312 22600 20343
rect 23382 20340 23388 20392
rect 23440 20380 23446 20392
rect 23477 20383 23535 20389
rect 23477 20380 23489 20383
rect 23440 20352 23489 20380
rect 23440 20340 23446 20352
rect 23477 20349 23489 20352
rect 23523 20349 23535 20383
rect 23477 20343 23535 20349
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20380 23811 20383
rect 24210 20380 24216 20392
rect 23799 20352 24216 20380
rect 23799 20349 23811 20352
rect 23753 20343 23811 20349
rect 24210 20340 24216 20352
rect 24268 20340 24274 20392
rect 20588 20284 21128 20312
rect 21192 20284 22600 20312
rect 20588 20272 20594 20284
rect 20070 20244 20076 20256
rect 18248 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 21192 20244 21220 20284
rect 20312 20216 21220 20244
rect 22005 20247 22063 20253
rect 20312 20204 20318 20216
rect 22005 20213 22017 20247
rect 22051 20244 22063 20247
rect 22370 20244 22376 20256
rect 22051 20216 22376 20244
rect 22051 20213 22063 20216
rect 22005 20207 22063 20213
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 25222 20204 25228 20256
rect 25280 20204 25286 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 6457 20043 6515 20049
rect 6457 20040 6469 20043
rect 4856 20012 6469 20040
rect 4856 20000 4862 20012
rect 6457 20009 6469 20012
rect 6503 20009 6515 20043
rect 6457 20003 6515 20009
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 7926 20040 7932 20052
rect 7064 20012 7932 20040
rect 7064 20000 7070 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10778 20040 10784 20052
rect 10192 20012 10784 20040
rect 10192 20000 10198 20012
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 11072 20012 14933 20040
rect 4982 19932 4988 19984
rect 5040 19972 5046 19984
rect 7101 19975 7159 19981
rect 7101 19972 7113 19975
rect 5040 19944 7113 19972
rect 5040 19932 5046 19944
rect 7101 19941 7113 19944
rect 7147 19941 7159 19975
rect 10594 19972 10600 19984
rect 7101 19935 7159 19941
rect 9324 19944 10600 19972
rect 2866 19864 2872 19916
rect 2924 19864 2930 19916
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19904 4859 19907
rect 5442 19904 5448 19916
rect 4847 19876 5448 19904
rect 4847 19873 4859 19876
rect 4801 19867 4859 19873
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 9324 19904 9352 19944
rect 10594 19932 10600 19944
rect 10652 19932 10658 19984
rect 6656 19876 9352 19904
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 3694 19836 3700 19848
rect 2271 19808 3700 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19836 4583 19839
rect 5902 19836 5908 19848
rect 4571 19808 5908 19836
rect 4571 19805 4583 19808
rect 4525 19799 4583 19805
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 6656 19845 6684 19876
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9769 19907 9827 19913
rect 9769 19904 9781 19907
rect 9456 19876 9781 19904
rect 9456 19864 9462 19876
rect 9769 19873 9781 19876
rect 9815 19904 9827 19907
rect 10870 19904 10876 19916
rect 9815 19876 10876 19904
rect 9815 19873 9827 19876
rect 9769 19867 9827 19873
rect 10870 19864 10876 19876
rect 10928 19864 10934 19916
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7466 19836 7472 19848
rect 7331 19808 7472 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 6012 19768 6040 19799
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7926 19796 7932 19848
rect 7984 19796 7990 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 9585 19839 9643 19845
rect 9585 19836 9597 19839
rect 8619 19808 9597 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 9585 19805 9597 19808
rect 9631 19805 9643 19839
rect 9585 19799 9643 19805
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19836 9735 19839
rect 11072 19836 11100 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 15010 20000 15016 20052
rect 15068 20040 15074 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 15068 20012 17693 20040
rect 15068 20000 15074 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 17770 20000 17776 20052
rect 17828 20040 17834 20052
rect 20254 20040 20260 20052
rect 17828 20012 20260 20040
rect 17828 20000 17834 20012
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 25038 20040 25044 20052
rect 21192 20012 25044 20040
rect 13354 19932 13360 19984
rect 13412 19932 13418 19984
rect 13722 19932 13728 19984
rect 13780 19972 13786 19984
rect 16301 19975 16359 19981
rect 16301 19972 16313 19975
rect 13780 19944 16313 19972
rect 13780 19932 13786 19944
rect 16301 19941 16313 19944
rect 16347 19941 16359 19975
rect 16301 19935 16359 19941
rect 16408 19944 18276 19972
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 13538 19904 13544 19916
rect 11655 19876 13544 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 13538 19864 13544 19876
rect 13596 19904 13602 19916
rect 14274 19904 14280 19916
rect 13596 19876 14280 19904
rect 13596 19864 13602 19876
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 14366 19864 14372 19916
rect 14424 19904 14430 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 14424 19876 15485 19904
rect 14424 19864 14430 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 16408 19904 16436 19944
rect 18248 19913 18276 19944
rect 18322 19932 18328 19984
rect 18380 19972 18386 19984
rect 21192 19972 21220 20012
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 18380 19944 21220 19972
rect 18380 19932 18386 19944
rect 22830 19932 22836 19984
rect 22888 19932 22894 19984
rect 15712 19876 16436 19904
rect 16853 19907 16911 19913
rect 15712 19864 15718 19876
rect 16853 19873 16865 19907
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19873 18291 19907
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 18233 19867 18291 19873
rect 18340 19876 19993 19904
rect 13630 19836 13636 19848
rect 9723 19808 11100 19836
rect 13372 19808 13636 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 13372 19780 13400 19808
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 13964 19808 14473 19836
rect 13964 19796 13970 19808
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 16868 19836 16896 19867
rect 14608 19808 16896 19836
rect 14608 19796 14614 19808
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 18340 19836 18368 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 22094 19904 22100 19916
rect 21131 19876 22100 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 22646 19864 22652 19916
rect 22704 19864 22710 19916
rect 25130 19864 25136 19916
rect 25188 19864 25194 19916
rect 18012 19808 18368 19836
rect 18012 19796 18018 19808
rect 19794 19796 19800 19848
rect 19852 19796 19858 19848
rect 22664 19836 22692 19864
rect 24302 19836 24308 19848
rect 22494 19822 24308 19836
rect 22480 19808 24308 19822
rect 6012 19740 9260 19768
rect 5813 19703 5871 19709
rect 5813 19669 5825 19703
rect 5859 19700 5871 19703
rect 6086 19700 6092 19712
rect 5859 19672 6092 19700
rect 5859 19669 5871 19672
rect 5813 19663 5871 19669
rect 6086 19660 6092 19672
rect 6144 19660 6150 19712
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 9232 19709 9260 19740
rect 9766 19728 9772 19780
rect 9824 19768 9830 19780
rect 11054 19768 11060 19780
rect 9824 19740 11060 19768
rect 9824 19728 9830 19740
rect 11054 19728 11060 19740
rect 11112 19728 11118 19780
rect 11882 19728 11888 19780
rect 11940 19728 11946 19780
rect 13354 19768 13360 19780
rect 13110 19740 13360 19768
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 13446 19728 13452 19780
rect 13504 19768 13510 19780
rect 15289 19771 15347 19777
rect 15289 19768 15301 19771
rect 13504 19740 15301 19768
rect 13504 19728 13510 19740
rect 15289 19737 15301 19740
rect 15335 19737 15347 19771
rect 15289 19731 15347 19737
rect 15378 19728 15384 19780
rect 15436 19728 15442 19780
rect 16669 19771 16727 19777
rect 16669 19737 16681 19771
rect 16715 19768 16727 19771
rect 17494 19768 17500 19780
rect 16715 19740 17500 19768
rect 16715 19737 16727 19740
rect 16669 19731 16727 19737
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 17586 19728 17592 19780
rect 17644 19768 17650 19780
rect 17880 19768 17908 19796
rect 18141 19771 18199 19777
rect 18141 19768 18153 19771
rect 17644 19740 18153 19768
rect 17644 19728 17650 19740
rect 18141 19737 18153 19740
rect 18187 19768 18199 19771
rect 19702 19768 19708 19780
rect 18187 19740 19708 19768
rect 18187 19737 18199 19740
rect 18141 19731 18199 19737
rect 19702 19728 19708 19740
rect 19760 19728 19766 19780
rect 21358 19728 21364 19780
rect 21416 19728 21422 19780
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7248 19672 7757 19700
rect 7248 19660 7254 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 9217 19703 9275 19709
rect 9217 19669 9229 19703
rect 9263 19669 9275 19703
rect 9217 19663 9275 19669
rect 10410 19660 10416 19712
rect 10468 19660 10474 19712
rect 10778 19660 10784 19712
rect 10836 19660 10842 19712
rect 10873 19703 10931 19709
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 12066 19700 12072 19712
rect 10919 19672 12072 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 12066 19660 12072 19672
rect 12124 19660 12130 19712
rect 14277 19703 14335 19709
rect 14277 19669 14289 19703
rect 14323 19700 14335 19703
rect 14366 19700 14372 19712
rect 14323 19672 14372 19700
rect 14323 19669 14335 19672
rect 14277 19663 14335 19669
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16298 19700 16304 19712
rect 16080 19672 16304 19700
rect 16080 19660 16086 19672
rect 16298 19660 16304 19672
rect 16356 19700 16362 19712
rect 16761 19703 16819 19709
rect 16761 19700 16773 19703
rect 16356 19672 16773 19700
rect 16356 19660 16362 19672
rect 16761 19669 16773 19672
rect 16807 19669 16819 19703
rect 16761 19663 16819 19669
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 18012 19672 18061 19700
rect 18012 19660 18018 19672
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18049 19663 18107 19669
rect 19426 19660 19432 19712
rect 19484 19660 19490 19712
rect 19889 19703 19947 19709
rect 19889 19669 19901 19703
rect 19935 19700 19947 19703
rect 19978 19700 19984 19712
rect 19935 19672 19984 19700
rect 19935 19669 19947 19672
rect 19889 19663 19947 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 22480 19700 22508 19808
rect 24302 19796 24308 19808
rect 24360 19796 24366 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19836 25007 19839
rect 25314 19836 25320 19848
rect 24995 19808 25320 19836
rect 24995 19805 25007 19808
rect 24949 19799 25007 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 25041 19771 25099 19777
rect 25041 19768 25053 19771
rect 23768 19740 25053 19768
rect 21140 19672 22508 19700
rect 21140 19660 21146 19672
rect 23290 19660 23296 19712
rect 23348 19700 23354 19712
rect 23768 19709 23796 19740
rect 25041 19737 25053 19740
rect 25087 19737 25099 19771
rect 25041 19731 25099 19737
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23348 19672 23765 19700
rect 23348 19660 23354 19672
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 24486 19660 24492 19712
rect 24544 19700 24550 19712
rect 24581 19703 24639 19709
rect 24581 19700 24593 19703
rect 24544 19672 24593 19700
rect 24544 19660 24550 19672
rect 24581 19669 24593 19672
rect 24627 19669 24639 19703
rect 24581 19663 24639 19669
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 3878 19456 3884 19508
rect 3936 19496 3942 19508
rect 4157 19499 4215 19505
rect 4157 19496 4169 19499
rect 3936 19468 4169 19496
rect 3936 19456 3942 19468
rect 4157 19465 4169 19468
rect 4203 19465 4215 19499
rect 4157 19459 4215 19465
rect 5442 19456 5448 19508
rect 5500 19456 5506 19508
rect 6178 19496 6184 19508
rect 6012 19468 6184 19496
rect 4798 19428 4804 19440
rect 4356 19400 4804 19428
rect 1946 19320 1952 19372
rect 2004 19320 2010 19372
rect 4356 19369 4384 19400
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19329 4399 19363
rect 4341 19323 4399 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 4764 19332 5580 19360
rect 4764 19320 4770 19332
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1728 19264 2237 19292
rect 1728 19252 1734 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 5552 19292 5580 19332
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 6012 19369 6040 19468
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 6549 19499 6607 19505
rect 6549 19465 6561 19499
rect 6595 19496 6607 19499
rect 7282 19496 7288 19508
rect 6595 19468 7288 19496
rect 6595 19465 6607 19468
rect 6549 19459 6607 19465
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 7742 19456 7748 19508
rect 7800 19456 7806 19508
rect 10410 19496 10416 19508
rect 7852 19468 10416 19496
rect 6638 19388 6644 19440
rect 6696 19428 6702 19440
rect 7852 19428 7880 19468
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 10870 19456 10876 19508
rect 10928 19456 10934 19508
rect 11882 19456 11888 19508
rect 11940 19496 11946 19508
rect 14461 19499 14519 19505
rect 14461 19496 14473 19499
rect 11940 19468 14473 19496
rect 11940 19456 11946 19468
rect 14461 19465 14473 19468
rect 14507 19496 14519 19499
rect 14550 19496 14556 19508
rect 14507 19468 14556 19496
rect 14507 19465 14519 19468
rect 14461 19459 14519 19465
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14884 19468 14933 19496
rect 14884 19456 14890 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 19426 19496 19432 19508
rect 15335 19468 16068 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 8478 19428 8484 19440
rect 6696 19400 7144 19428
rect 6696 19388 6702 19400
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19329 6055 19363
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 5997 19323 6055 19329
rect 6104 19332 6745 19360
rect 6104 19292 6132 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 5552 19264 6132 19292
rect 2225 19255 2283 19261
rect 5353 19227 5411 19233
rect 5353 19193 5365 19227
rect 5399 19224 5411 19227
rect 6178 19224 6184 19236
rect 5399 19196 6184 19224
rect 5399 19193 5411 19196
rect 5353 19187 5411 19193
rect 6178 19184 6184 19196
rect 6236 19184 6242 19236
rect 4065 19159 4123 19165
rect 4065 19125 4077 19159
rect 4111 19156 4123 19159
rect 4706 19156 4712 19168
rect 4111 19128 4712 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5813 19159 5871 19165
rect 5813 19125 5825 19159
rect 5859 19156 5871 19159
rect 6270 19156 6276 19168
rect 5859 19128 6276 19156
rect 5859 19125 5871 19128
rect 5813 19119 5871 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 7116 19156 7144 19400
rect 7392 19400 7880 19428
rect 7944 19400 8484 19428
rect 7392 19369 7420 19400
rect 7944 19369 7972 19400
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 11514 19388 11520 19440
rect 11572 19428 11578 19440
rect 13262 19428 13268 19440
rect 11572 19400 13268 19428
rect 11572 19388 11578 19400
rect 13262 19388 13268 19400
rect 13320 19388 13326 19440
rect 13446 19388 13452 19440
rect 13504 19388 13510 19440
rect 15010 19388 15016 19440
rect 15068 19428 15074 19440
rect 15654 19428 15660 19440
rect 15068 19400 15660 19428
rect 15068 19388 15074 19400
rect 15654 19388 15660 19400
rect 15712 19388 15718 19440
rect 16040 19428 16068 19468
rect 16316 19468 19432 19496
rect 16316 19428 16344 19468
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 20349 19499 20407 19505
rect 20349 19465 20361 19499
rect 20395 19496 20407 19499
rect 20714 19496 20720 19508
rect 20395 19468 20720 19496
rect 20395 19465 20407 19468
rect 20349 19459 20407 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 22005 19499 22063 19505
rect 22005 19465 22017 19499
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 16574 19428 16580 19440
rect 16040 19400 16344 19428
rect 16408 19400 16580 19428
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19329 8263 19363
rect 8205 19323 8263 19329
rect 8018 19292 8024 19304
rect 7208 19264 8024 19292
rect 7208 19233 7236 19264
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 8220 19292 8248 19323
rect 10502 19320 10508 19372
rect 10560 19320 10566 19372
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 12069 19363 12127 19369
rect 12069 19360 12081 19363
rect 11756 19332 12081 19360
rect 11756 19320 11762 19332
rect 12069 19329 12081 19332
rect 12115 19329 12127 19363
rect 12069 19323 12127 19329
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12710 19360 12716 19372
rect 12400 19332 12716 19360
rect 12400 19320 12406 19332
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 16264 19332 16313 19360
rect 16264 19320 16270 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 8478 19292 8484 19304
rect 8220 19264 8484 19292
rect 8478 19252 8484 19264
rect 8536 19252 8542 19304
rect 9122 19252 9128 19304
rect 9180 19252 9186 19304
rect 9401 19295 9459 19301
rect 9401 19261 9413 19295
rect 9447 19292 9459 19295
rect 10686 19292 10692 19304
rect 9447 19264 10692 19292
rect 9447 19261 9459 19264
rect 9401 19255 9459 19261
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 15102 19292 15108 19304
rect 13035 19264 15108 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15378 19252 15384 19304
rect 15436 19252 15442 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16022 19292 16028 19304
rect 15611 19264 16028 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 7193 19227 7251 19233
rect 7193 19193 7205 19227
rect 7239 19193 7251 19227
rect 7193 19187 7251 19193
rect 10410 19184 10416 19236
rect 10468 19224 10474 19236
rect 10468 19196 10903 19224
rect 10468 19184 10474 19196
rect 8021 19159 8079 19165
rect 8021 19156 8033 19159
rect 7116 19128 8033 19156
rect 8021 19125 8033 19128
rect 8067 19125 8079 19159
rect 8021 19119 8079 19125
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19156 8723 19159
rect 10778 19156 10784 19168
rect 8711 19128 10784 19156
rect 8711 19125 8723 19128
rect 8665 19119 8723 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 10875 19156 10903 19196
rect 11054 19184 11060 19236
rect 11112 19224 11118 19236
rect 16408 19224 16436 19400
rect 16574 19388 16580 19400
rect 16632 19388 16638 19440
rect 17954 19388 17960 19440
rect 18012 19388 18018 19440
rect 19521 19431 19579 19437
rect 19521 19397 19533 19431
rect 19567 19428 19579 19431
rect 20530 19428 20536 19440
rect 19567 19400 20536 19428
rect 19567 19397 19579 19400
rect 19521 19391 19579 19397
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 22020 19428 22048 19459
rect 22370 19456 22376 19508
rect 22428 19456 22434 19508
rect 22465 19499 22523 19505
rect 22465 19465 22477 19499
rect 22511 19496 22523 19499
rect 22554 19496 22560 19508
rect 22511 19468 22560 19496
rect 22511 19465 22523 19468
rect 22465 19459 22523 19465
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 25133 19499 25191 19505
rect 25133 19465 25145 19499
rect 25179 19496 25191 19499
rect 25406 19496 25412 19508
rect 25179 19468 25412 19496
rect 25179 19465 25191 19468
rect 25133 19459 25191 19465
rect 25406 19456 25412 19468
rect 25464 19456 25470 19508
rect 23658 19428 23664 19440
rect 22020 19400 23664 19428
rect 23658 19388 23664 19400
rect 23716 19388 23722 19440
rect 24302 19388 24308 19440
rect 24360 19388 24366 19440
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 16945 19363 17003 19369
rect 16945 19360 16957 19363
rect 16540 19332 16957 19360
rect 16540 19320 16546 19332
rect 16945 19329 16957 19332
rect 16991 19329 17003 19363
rect 19426 19360 19432 19372
rect 16945 19323 17003 19329
rect 18708 19332 19432 19360
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 16632 19264 17233 19292
rect 16632 19252 16638 19264
rect 17221 19261 17233 19264
rect 17267 19292 17279 19295
rect 17678 19292 17684 19304
rect 17267 19264 17684 19292
rect 17267 19261 17279 19264
rect 17221 19255 17279 19261
rect 17678 19252 17684 19264
rect 17736 19252 17742 19304
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18506 19292 18512 19304
rect 18012 19264 18512 19292
rect 18012 19252 18018 19264
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 18708 19301 18736 19332
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 20622 19320 20628 19372
rect 20680 19360 20686 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20680 19332 20729 19360
rect 20680 19320 20686 19332
rect 20717 19329 20729 19332
rect 20763 19360 20775 19363
rect 21818 19360 21824 19372
rect 20763 19332 21824 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19261 18751 19295
rect 19444 19292 19472 19320
rect 19444 19264 19564 19292
rect 18693 19255 18751 19261
rect 19334 19224 19340 19236
rect 11112 19196 12296 19224
rect 11112 19184 11118 19196
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 10875 19128 12173 19156
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 12268 19156 12296 19196
rect 16224 19196 16436 19224
rect 18248 19196 19340 19224
rect 13446 19156 13452 19168
rect 12268 19128 13452 19156
rect 12161 19119 12219 19125
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 15286 19156 15292 19168
rect 14608 19128 15292 19156
rect 14608 19116 14614 19128
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16224 19156 16252 19196
rect 16163 19128 16252 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 17034 19116 17040 19168
rect 17092 19156 17098 19168
rect 18248 19156 18276 19196
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 19536 19224 19564 19264
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19292 21051 19295
rect 22002 19292 22008 19304
rect 21039 19264 22008 19292
rect 21039 19261 21051 19264
rect 20993 19255 21051 19261
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 22572 19224 22600 19255
rect 23382 19252 23388 19304
rect 23440 19252 23446 19304
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 25222 19292 25228 19304
rect 23707 19264 25228 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 19536 19196 22600 19224
rect 17092 19128 18276 19156
rect 19153 19159 19211 19165
rect 17092 19116 17098 19128
rect 19153 19125 19165 19159
rect 19199 19156 19211 19159
rect 19518 19156 19524 19168
rect 19199 19128 19524 19156
rect 19199 19125 19211 19128
rect 19153 19119 19211 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21174 19156 21180 19168
rect 20956 19128 21180 19156
rect 20956 19116 20962 19128
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 22520 19128 23213 19156
rect 22520 19116 22526 19128
rect 23201 19125 23213 19128
rect 23247 19156 23259 19159
rect 24762 19156 24768 19168
rect 23247 19128 24768 19156
rect 23247 19125 23259 19128
rect 23201 19119 23259 19125
rect 24762 19116 24768 19128
rect 24820 19116 24826 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 1949 18955 2007 18961
rect 1949 18921 1961 18955
rect 1995 18952 2007 18955
rect 2130 18952 2136 18964
rect 1995 18924 2136 18952
rect 1995 18921 2007 18924
rect 1949 18915 2007 18921
rect 2130 18912 2136 18924
rect 2188 18912 2194 18964
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 14277 18955 14335 18961
rect 4764 18924 14228 18952
rect 4764 18912 4770 18924
rect 4522 18844 4528 18896
rect 4580 18884 4586 18896
rect 5445 18887 5503 18893
rect 5445 18884 5457 18887
rect 4580 18856 5457 18884
rect 4580 18844 4586 18856
rect 5445 18853 5457 18856
rect 5491 18853 5503 18887
rect 5445 18847 5503 18853
rect 5626 18844 5632 18896
rect 5684 18884 5690 18896
rect 5813 18887 5871 18893
rect 5813 18884 5825 18887
rect 5684 18856 5825 18884
rect 5684 18844 5690 18856
rect 5813 18853 5825 18856
rect 5859 18853 5871 18887
rect 8386 18884 8392 18896
rect 5813 18847 5871 18853
rect 5920 18856 8392 18884
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18816 4307 18819
rect 5350 18816 5356 18828
rect 4295 18788 5356 18816
rect 4295 18785 4307 18788
rect 4249 18779 4307 18785
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 2133 18751 2191 18757
rect 2133 18748 2145 18751
rect 1903 18720 2145 18748
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 2133 18717 2145 18720
rect 2179 18748 2191 18751
rect 2222 18748 2228 18760
rect 2179 18720 2228 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18748 2927 18751
rect 3513 18751 3571 18757
rect 3513 18748 3525 18751
rect 2915 18720 3525 18748
rect 2915 18717 2927 18720
rect 2869 18711 2927 18717
rect 3513 18717 3525 18720
rect 3559 18748 3571 18751
rect 4338 18748 4344 18760
rect 3559 18720 4344 18748
rect 3559 18717 3571 18720
rect 3513 18711 3571 18717
rect 4338 18708 4344 18720
rect 4396 18708 4402 18760
rect 4724 18757 4752 18788
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18748 5687 18751
rect 5920 18748 5948 18856
rect 8386 18844 8392 18856
rect 8444 18844 8450 18896
rect 8846 18884 8852 18896
rect 8496 18856 8852 18884
rect 7834 18816 7840 18828
rect 6012 18788 7840 18816
rect 6012 18757 6040 18788
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 8496 18816 8524 18856
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 14200 18884 14228 18924
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 15378 18952 15384 18964
rect 14323 18924 15384 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 15488 18924 16804 18952
rect 15488 18884 15516 18924
rect 14200 18856 15516 18884
rect 16776 18884 16804 18924
rect 17218 18912 17224 18964
rect 17276 18912 17282 18964
rect 18782 18912 18788 18964
rect 18840 18952 18846 18964
rect 19702 18952 19708 18964
rect 18840 18924 19708 18952
rect 18840 18912 18846 18924
rect 19702 18912 19708 18924
rect 19760 18912 19766 18964
rect 19812 18924 23060 18952
rect 18414 18884 18420 18896
rect 16776 18856 18420 18884
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 18874 18844 18880 18896
rect 18932 18884 18938 18896
rect 19812 18884 19840 18924
rect 18932 18856 19840 18884
rect 18932 18844 18938 18856
rect 7984 18788 8524 18816
rect 8665 18819 8723 18825
rect 7984 18776 7990 18788
rect 8665 18785 8677 18819
rect 8711 18816 8723 18819
rect 8711 18788 11100 18816
rect 8711 18785 8723 18788
rect 8665 18779 8723 18785
rect 5675 18720 5948 18748
rect 5997 18751 6055 18757
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 5997 18717 6009 18751
rect 6043 18717 6055 18751
rect 5997 18711 6055 18717
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 7285 18751 7343 18757
rect 7285 18717 7297 18751
rect 7331 18748 7343 18751
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7331 18720 8401 18748
rect 7331 18717 7343 18720
rect 7285 18711 7343 18717
rect 8389 18717 8401 18720
rect 8435 18748 8447 18751
rect 8754 18748 8760 18760
rect 8435 18720 8760 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 10502 18708 10508 18760
rect 10560 18708 10566 18760
rect 11072 18748 11100 18788
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 11204 18788 11713 18816
rect 11204 18776 11210 18788
rect 11701 18785 11713 18788
rect 11747 18816 11759 18819
rect 11974 18816 11980 18828
rect 11747 18788 11980 18816
rect 11747 18785 11759 18788
rect 11701 18779 11759 18785
rect 11974 18776 11980 18788
rect 12032 18816 12038 18828
rect 12342 18816 12348 18828
rect 12032 18788 12348 18816
rect 12032 18776 12038 18788
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 13446 18816 13452 18828
rect 12584 18788 13452 18816
rect 12584 18776 12590 18788
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14918 18816 14924 18828
rect 14148 18788 14924 18816
rect 14148 18776 14154 18788
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 16482 18816 16488 18828
rect 15488 18788 16488 18816
rect 11606 18748 11612 18760
rect 11072 18720 11612 18748
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 14274 18708 14280 18760
rect 14332 18748 14338 18760
rect 15488 18757 15516 18788
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 18322 18776 18328 18828
rect 18380 18776 18386 18828
rect 19242 18776 19248 18828
rect 19300 18816 19306 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 19300 18788 20361 18816
rect 19300 18776 19306 18788
rect 20349 18785 20361 18788
rect 20395 18785 20407 18819
rect 20349 18779 20407 18785
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18816 20683 18819
rect 22830 18816 22836 18828
rect 20671 18788 22836 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 23032 18825 23060 18924
rect 23385 18887 23443 18893
rect 23124 18856 23336 18884
rect 23017 18819 23075 18825
rect 23017 18785 23029 18819
rect 23063 18785 23075 18819
rect 23017 18779 23075 18785
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 14332 18720 15485 18748
rect 14332 18708 14338 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 18046 18708 18052 18760
rect 18104 18708 18110 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19886 18748 19892 18760
rect 19659 18720 19892 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 22554 18708 22560 18760
rect 22612 18748 22618 18760
rect 23124 18748 23152 18856
rect 23201 18819 23259 18825
rect 23201 18785 23213 18819
rect 23247 18785 23259 18819
rect 23201 18779 23259 18785
rect 22612 18720 23152 18748
rect 22612 18708 22618 18720
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18680 5411 18683
rect 6656 18680 6684 18708
rect 8202 18680 8208 18692
rect 5399 18652 6684 18680
rect 7024 18652 8208 18680
rect 5399 18649 5411 18652
rect 5353 18643 5411 18649
rect 3329 18615 3387 18621
rect 3329 18581 3341 18615
rect 3375 18612 3387 18615
rect 4062 18612 4068 18624
rect 3375 18584 4068 18612
rect 3375 18581 3387 18584
rect 3329 18575 3387 18581
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 4525 18615 4583 18621
rect 4525 18581 4537 18615
rect 4571 18612 4583 18615
rect 7024 18612 7052 18652
rect 8202 18640 8208 18652
rect 8260 18640 8266 18692
rect 9398 18640 9404 18692
rect 9456 18640 9462 18692
rect 11238 18680 11244 18692
rect 9508 18652 9812 18680
rect 9508 18624 9536 18652
rect 4571 18584 7052 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 7098 18572 7104 18624
rect 7156 18572 7162 18624
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 9122 18612 9128 18624
rect 7340 18584 9128 18612
rect 7340 18572 7346 18584
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 9490 18572 9496 18624
rect 9548 18572 9554 18624
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 9674 18612 9680 18624
rect 9640 18584 9680 18612
rect 9640 18572 9646 18584
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 9784 18612 9812 18652
rect 10704 18652 11244 18680
rect 10704 18612 10732 18652
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 11514 18640 11520 18692
rect 11572 18680 11578 18692
rect 11977 18683 12035 18689
rect 11977 18680 11989 18683
rect 11572 18652 11989 18680
rect 11572 18640 11578 18652
rect 11977 18649 11989 18652
rect 12023 18680 12035 18683
rect 12250 18680 12256 18692
rect 12023 18652 12256 18680
rect 12023 18649 12035 18652
rect 11977 18643 12035 18649
rect 12250 18640 12256 18652
rect 12308 18640 12314 18692
rect 12710 18640 12716 18692
rect 12768 18640 12774 18692
rect 15749 18683 15807 18689
rect 13372 18652 14872 18680
rect 9784 18584 10732 18612
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 13372 18612 13400 18652
rect 10928 18584 13400 18612
rect 10928 18572 10934 18584
rect 13446 18572 13452 18624
rect 13504 18572 13510 18624
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 14608 18584 14657 18612
rect 14608 18572 14614 18584
rect 14645 18581 14657 18584
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 14734 18572 14740 18624
rect 14792 18572 14798 18624
rect 14844 18612 14872 18652
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16022 18680 16028 18692
rect 15795 18652 16028 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16206 18680 16212 18692
rect 16132 18652 16212 18680
rect 15838 18612 15844 18624
rect 14844 18584 15844 18612
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16132 18612 16160 18652
rect 16206 18640 16212 18652
rect 16264 18640 16270 18692
rect 17954 18680 17960 18692
rect 17604 18652 17960 18680
rect 17604 18612 17632 18652
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 21082 18640 21088 18692
rect 21140 18640 21146 18692
rect 23216 18680 23244 18779
rect 23308 18748 23336 18856
rect 23385 18853 23397 18887
rect 23431 18884 23443 18887
rect 24854 18884 24860 18896
rect 23431 18856 24860 18884
rect 23431 18853 23443 18856
rect 23385 18847 23443 18853
rect 24854 18844 24860 18856
rect 24912 18844 24918 18896
rect 23842 18776 23848 18828
rect 23900 18776 23906 18828
rect 24026 18776 24032 18828
rect 24084 18776 24090 18828
rect 25222 18776 25228 18828
rect 25280 18776 25286 18828
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23308 18720 23765 18748
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 24762 18708 24768 18760
rect 24820 18748 24826 18760
rect 24949 18751 25007 18757
rect 24949 18748 24961 18751
rect 24820 18720 24961 18748
rect 24820 18708 24826 18720
rect 24949 18717 24961 18720
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 25314 18680 25320 18692
rect 21928 18652 23244 18680
rect 23676 18652 25320 18680
rect 16132 18584 17632 18612
rect 17678 18572 17684 18624
rect 17736 18572 17742 18624
rect 18141 18615 18199 18621
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 19429 18615 19487 18621
rect 19429 18612 19441 18615
rect 18187 18584 19441 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 19429 18581 19441 18584
rect 19475 18581 19487 18615
rect 19429 18575 19487 18581
rect 20162 18572 20168 18624
rect 20220 18612 20226 18624
rect 21928 18612 21956 18652
rect 20220 18584 21956 18612
rect 22097 18615 22155 18621
rect 20220 18572 20226 18584
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22278 18612 22284 18624
rect 22143 18584 22284 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22554 18572 22560 18624
rect 22612 18572 22618 18624
rect 22922 18572 22928 18624
rect 22980 18612 22986 18624
rect 23676 18612 23704 18652
rect 25314 18640 25320 18652
rect 25372 18640 25378 18692
rect 22980 18584 23704 18612
rect 22980 18572 22986 18584
rect 24118 18572 24124 18624
rect 24176 18612 24182 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 24176 18584 24593 18612
rect 24176 18572 24182 18584
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 25038 18572 25044 18624
rect 25096 18572 25102 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 1857 18411 1915 18417
rect 1857 18377 1869 18411
rect 1903 18408 1915 18411
rect 6822 18408 6828 18420
rect 1903 18380 6828 18408
rect 1903 18377 1915 18380
rect 1857 18371 1915 18377
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 7374 18368 7380 18420
rect 7432 18408 7438 18420
rect 8021 18411 8079 18417
rect 8021 18408 8033 18411
rect 7432 18380 8033 18408
rect 7432 18368 7438 18380
rect 8021 18377 8033 18380
rect 8067 18377 8079 18411
rect 8021 18371 8079 18377
rect 8389 18411 8447 18417
rect 8389 18377 8401 18411
rect 8435 18408 8447 18411
rect 9030 18408 9036 18420
rect 8435 18380 9036 18408
rect 8435 18377 8447 18380
rect 8389 18371 8447 18377
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9122 18368 9128 18420
rect 9180 18368 9186 18420
rect 9600 18380 13032 18408
rect 4709 18343 4767 18349
rect 4709 18309 4721 18343
rect 4755 18340 4767 18343
rect 8846 18340 8852 18352
rect 4755 18312 5304 18340
rect 4755 18309 4767 18312
rect 4709 18303 4767 18309
rect 5276 18284 5304 18312
rect 8496 18312 8852 18340
rect 2038 18232 2044 18284
rect 2096 18232 2102 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 3326 18272 3332 18284
rect 2179 18244 3332 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18272 3571 18275
rect 4157 18275 4215 18281
rect 4157 18272 4169 18275
rect 3559 18244 4169 18272
rect 3559 18241 3571 18244
rect 3513 18235 3571 18241
rect 4157 18241 4169 18244
rect 4203 18272 4215 18275
rect 4430 18272 4436 18284
rect 4203 18244 4436 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4430 18232 4436 18244
rect 4488 18232 4494 18284
rect 4890 18272 4896 18284
rect 4540 18244 4896 18272
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 4540 18204 4568 18244
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 4982 18232 4988 18284
rect 5040 18232 5046 18284
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5353 18275 5411 18281
rect 5353 18272 5365 18275
rect 5316 18244 5365 18272
rect 5316 18232 5322 18244
rect 5353 18241 5365 18244
rect 5399 18241 5411 18275
rect 5353 18235 5411 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 7190 18272 7196 18284
rect 6043 18244 7196 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 7282 18232 7288 18284
rect 7340 18232 7346 18284
rect 8213 18275 8271 18281
rect 8213 18241 8225 18275
rect 8259 18272 8271 18275
rect 8496 18272 8524 18312
rect 8846 18300 8852 18312
rect 8904 18300 8910 18352
rect 9600 18284 9628 18380
rect 11146 18300 11152 18352
rect 11204 18300 11210 18352
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 12161 18343 12219 18349
rect 12161 18340 12173 18343
rect 11664 18312 12173 18340
rect 11664 18300 11670 18312
rect 12161 18309 12173 18312
rect 12207 18309 12219 18343
rect 12161 18303 12219 18309
rect 12250 18300 12256 18352
rect 12308 18340 12314 18352
rect 13004 18349 13032 18380
rect 14274 18368 14280 18420
rect 14332 18368 14338 18420
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17310 18408 17316 18420
rect 17267 18380 17316 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 19242 18408 19248 18420
rect 18472 18380 19248 18408
rect 18472 18368 18478 18380
rect 19242 18368 19248 18380
rect 19300 18408 19306 18420
rect 19521 18411 19579 18417
rect 19521 18408 19533 18411
rect 19300 18380 19533 18408
rect 19300 18368 19306 18380
rect 19521 18377 19533 18380
rect 19567 18377 19579 18411
rect 19521 18371 19579 18377
rect 20809 18411 20867 18417
rect 20809 18377 20821 18411
rect 20855 18408 20867 18411
rect 20898 18408 20904 18420
rect 20855 18380 20904 18408
rect 20855 18377 20867 18380
rect 20809 18371 20867 18377
rect 20898 18368 20904 18380
rect 20956 18408 20962 18420
rect 20956 18380 22692 18408
rect 20956 18368 20962 18380
rect 12989 18343 13047 18349
rect 12308 18312 12664 18340
rect 12308 18300 12314 18312
rect 8259 18244 8524 18272
rect 8573 18275 8631 18281
rect 8259 18241 8271 18244
rect 8213 18235 8271 18241
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8662 18272 8668 18284
rect 8619 18244 8668 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18272 9459 18275
rect 9582 18272 9588 18284
rect 9447 18244 9588 18272
rect 9447 18241 9459 18244
rect 9401 18235 9459 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 11422 18272 11428 18284
rect 10008 18244 11428 18272
rect 10008 18232 10014 18244
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 12526 18272 12532 18284
rect 12268 18244 12532 18272
rect 2455 18176 4568 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 4614 18164 4620 18216
rect 4672 18204 4678 18216
rect 4672 18176 4844 18204
rect 4672 18164 4678 18176
rect 3973 18139 4031 18145
rect 3973 18105 3985 18139
rect 4019 18136 4031 18139
rect 4706 18136 4712 18148
rect 4019 18108 4712 18136
rect 4019 18105 4031 18108
rect 3973 18099 4031 18105
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 4816 18145 4844 18176
rect 7926 18164 7932 18216
rect 7984 18164 7990 18216
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 10778 18204 10784 18216
rect 8444 18176 10784 18204
rect 8444 18164 8450 18176
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 12268 18213 12296 18244
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 12636 18272 12664 18312
rect 12989 18309 13001 18343
rect 13035 18340 13047 18343
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 13035 18312 18245 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 18233 18309 18245 18312
rect 18279 18340 18291 18343
rect 18506 18340 18512 18352
rect 18279 18312 18512 18340
rect 18279 18309 18291 18312
rect 18233 18303 18291 18309
rect 18506 18300 18512 18312
rect 18564 18340 18570 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 18564 18312 22017 18340
rect 18564 18300 18570 18312
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22664 18340 22692 18380
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 24581 18411 24639 18417
rect 24581 18408 24593 18411
rect 22796 18380 24593 18408
rect 22796 18368 22802 18380
rect 24581 18377 24593 18380
rect 24627 18377 24639 18411
rect 24581 18371 24639 18377
rect 24946 18368 24952 18420
rect 25004 18368 25010 18420
rect 22922 18340 22928 18352
rect 22664 18312 22928 18340
rect 22005 18303 22063 18309
rect 22922 18300 22928 18312
rect 22980 18300 22986 18352
rect 25038 18340 25044 18352
rect 23584 18312 25044 18340
rect 15010 18272 15016 18284
rect 12636 18244 15016 18272
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 15562 18232 15568 18284
rect 15620 18232 15626 18284
rect 16298 18272 16304 18284
rect 15672 18244 16304 18272
rect 15672 18216 15700 18244
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17313 18275 17371 18281
rect 17313 18272 17325 18275
rect 17184 18244 17325 18272
rect 17184 18232 17190 18244
rect 17313 18241 17325 18244
rect 17359 18272 17371 18275
rect 19886 18272 19892 18284
rect 17359 18244 19892 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20898 18232 20904 18284
rect 20956 18232 20962 18284
rect 23584 18272 23612 18312
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 21008 18244 23612 18272
rect 24121 18275 24179 18281
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 14734 18164 14740 18216
rect 14792 18204 14798 18216
rect 15654 18204 15660 18216
rect 14792 18176 15660 18204
rect 14792 18164 14798 18176
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 15838 18164 15844 18216
rect 15896 18164 15902 18216
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 21008 18204 21036 18244
rect 24121 18241 24133 18275
rect 24167 18272 24179 18275
rect 24762 18272 24768 18284
rect 24167 18244 24768 18272
rect 24167 18241 24179 18244
rect 24121 18235 24179 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 20404 18176 21036 18204
rect 20404 18164 20410 18176
rect 21082 18164 21088 18216
rect 21140 18164 21146 18216
rect 22830 18164 22836 18216
rect 22888 18204 22894 18216
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 22888 18176 25053 18204
rect 22888 18164 22894 18176
rect 25041 18173 25053 18176
rect 25087 18173 25099 18207
rect 25041 18167 25099 18173
rect 25133 18207 25191 18213
rect 25133 18173 25145 18207
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 4801 18139 4859 18145
rect 4801 18105 4813 18139
rect 4847 18105 4859 18139
rect 4801 18099 4859 18105
rect 5166 18096 5172 18148
rect 5224 18096 5230 18148
rect 5718 18096 5724 18148
rect 5776 18136 5782 18148
rect 5813 18139 5871 18145
rect 5813 18136 5825 18139
rect 5776 18108 5825 18136
rect 5776 18096 5782 18108
rect 5813 18105 5825 18108
rect 5859 18105 5871 18139
rect 5813 18099 5871 18105
rect 6638 18096 6644 18148
rect 6696 18136 6702 18148
rect 11054 18136 11060 18148
rect 6696 18108 11060 18136
rect 6696 18096 6702 18108
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 12584 18108 16865 18136
rect 12584 18096 12590 18108
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 16853 18099 16911 18105
rect 17218 18096 17224 18148
rect 17276 18136 17282 18148
rect 23937 18139 23995 18145
rect 23937 18136 23949 18139
rect 17276 18108 23949 18136
rect 17276 18096 17282 18108
rect 23937 18105 23949 18108
rect 23983 18105 23995 18139
rect 23937 18099 23995 18105
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 6914 18068 6920 18080
rect 5408 18040 6920 18068
rect 5408 18028 5414 18040
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 7101 18071 7159 18077
rect 7101 18037 7113 18071
rect 7147 18068 7159 18071
rect 9398 18068 9404 18080
rect 7147 18040 9404 18068
rect 7147 18037 7159 18040
rect 7101 18031 7159 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 10652 18040 11805 18068
rect 10652 18028 10658 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12066 18028 12072 18080
rect 12124 18068 12130 18080
rect 15197 18071 15255 18077
rect 15197 18068 15209 18071
rect 12124 18040 15209 18068
rect 12124 18028 12130 18040
rect 15197 18037 15209 18040
rect 15243 18037 15255 18071
rect 15197 18031 15255 18037
rect 15562 18028 15568 18080
rect 15620 18068 15626 18080
rect 16206 18068 16212 18080
rect 15620 18040 16212 18068
rect 15620 18028 15626 18040
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 20622 18068 20628 18080
rect 20487 18040 20628 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 23293 18071 23351 18077
rect 23293 18068 23305 18071
rect 22152 18040 23305 18068
rect 22152 18028 22158 18040
rect 23293 18037 23305 18040
rect 23339 18068 23351 18071
rect 23382 18068 23388 18080
rect 23339 18040 23388 18068
rect 23339 18037 23351 18040
rect 23293 18031 23351 18037
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 25148 18068 25176 18167
rect 23624 18040 25176 18068
rect 23624 18028 23630 18040
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 2096 17836 2145 17864
rect 2096 17824 2102 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 2133 17827 2191 17833
rect 5074 17824 5080 17876
rect 5132 17864 5138 17876
rect 5169 17867 5227 17873
rect 5169 17864 5181 17867
rect 5132 17836 5181 17864
rect 5132 17824 5138 17836
rect 5169 17833 5181 17836
rect 5215 17833 5227 17867
rect 5169 17827 5227 17833
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 5592 17836 6745 17864
rect 5592 17824 5598 17836
rect 6733 17833 6745 17836
rect 6779 17833 6791 17867
rect 6733 17827 6791 17833
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7708 17836 7757 17864
rect 7708 17824 7714 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 7745 17827 7803 17833
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 15838 17864 15844 17876
rect 8435 17836 15844 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 15838 17824 15844 17836
rect 15896 17824 15902 17876
rect 16574 17824 16580 17876
rect 16632 17824 16638 17876
rect 18233 17867 18291 17873
rect 18233 17833 18245 17867
rect 18279 17864 18291 17867
rect 18690 17864 18696 17876
rect 18279 17836 18696 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18690 17824 18696 17836
rect 18748 17824 18754 17876
rect 21358 17824 21364 17876
rect 21416 17864 21422 17876
rect 21416 17836 21864 17864
rect 21416 17824 21422 17836
rect 7098 17756 7104 17808
rect 7156 17756 7162 17808
rect 9125 17799 9183 17805
rect 9125 17796 9137 17799
rect 7208 17768 9137 17796
rect 5994 17688 6000 17740
rect 6052 17728 6058 17740
rect 7208 17728 7236 17768
rect 9125 17765 9137 17768
rect 9171 17765 9183 17799
rect 9125 17759 9183 17765
rect 11514 17756 11520 17808
rect 11572 17756 11578 17808
rect 13722 17756 13728 17808
rect 13780 17796 13786 17808
rect 17402 17796 17408 17808
rect 13780 17768 14964 17796
rect 13780 17756 13786 17768
rect 6052 17700 7236 17728
rect 8588 17700 11652 17728
rect 6052 17688 6058 17700
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 3421 17663 3479 17669
rect 3421 17660 3433 17663
rect 2823 17632 3433 17660
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 3421 17629 3433 17632
rect 3467 17660 3479 17663
rect 3786 17660 3792 17672
rect 3467 17632 3792 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3786 17620 3792 17632
rect 3844 17620 3850 17672
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 5074 17660 5080 17672
rect 4755 17632 5080 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 5868 17632 6929 17660
rect 5868 17620 5874 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 3694 17552 3700 17604
rect 3752 17592 3758 17604
rect 6641 17595 6699 17601
rect 3752 17564 4660 17592
rect 3752 17552 3758 17564
rect 3234 17484 3240 17536
rect 3292 17484 3298 17536
rect 4522 17484 4528 17536
rect 4580 17484 4586 17536
rect 4632 17524 4660 17564
rect 6641 17561 6653 17595
rect 6687 17592 6699 17595
rect 7300 17592 7328 17623
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 8588 17669 8616 17700
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7800 17632 7941 17660
rect 7800 17620 7806 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 9309 17663 9367 17669
rect 9309 17660 9321 17663
rect 9272 17632 9321 17660
rect 9272 17620 9278 17632
rect 9309 17629 9321 17632
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9732 17632 9781 17660
rect 9732 17620 9738 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 11146 17620 11152 17672
rect 11204 17620 11210 17672
rect 8754 17592 8760 17604
rect 6687 17564 8760 17592
rect 6687 17561 6699 17564
rect 6641 17555 6699 17561
rect 8754 17552 8760 17564
rect 8812 17552 8818 17604
rect 10045 17595 10103 17601
rect 10045 17561 10057 17595
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 9858 17524 9864 17536
rect 4632 17496 9864 17524
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 10060 17524 10088 17555
rect 10962 17524 10968 17536
rect 10060 17496 10968 17524
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11624 17524 11652 17700
rect 11974 17688 11980 17740
rect 12032 17688 12038 17740
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12618 17728 12624 17740
rect 12299 17700 12624 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12618 17688 12624 17700
rect 12676 17728 12682 17740
rect 13446 17728 13452 17740
rect 12676 17700 13452 17728
rect 12676 17688 12682 17700
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14829 17731 14887 17737
rect 14829 17728 14841 17731
rect 14332 17700 14841 17728
rect 14332 17688 14338 17700
rect 14829 17697 14841 17700
rect 14875 17697 14887 17731
rect 14936 17728 14964 17768
rect 16132 17768 17408 17796
rect 16132 17728 16160 17768
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 21836 17796 21864 17836
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 23382 17864 23388 17876
rect 21968 17836 23388 17864
rect 21968 17824 21974 17836
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 21836 17768 23888 17796
rect 23860 17740 23888 17768
rect 14936 17700 16160 17728
rect 14829 17691 14887 17697
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 16632 17700 17601 17728
rect 16632 17688 16638 17700
rect 17589 17697 17601 17700
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 17696 17700 19380 17728
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 17696 17660 17724 17700
rect 16540 17632 17724 17660
rect 18417 17663 18475 17669
rect 16540 17620 16546 17632
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 19242 17660 19248 17672
rect 18463 17632 19248 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 19352 17660 19380 17700
rect 19610 17688 19616 17740
rect 19668 17728 19674 17740
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 19668 17700 19993 17728
rect 19668 17688 19674 17700
rect 19981 17697 19993 17700
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20533 17731 20591 17737
rect 20533 17697 20545 17731
rect 20579 17728 20591 17731
rect 22094 17728 22100 17740
rect 20579 17700 22100 17728
rect 20579 17697 20591 17700
rect 20533 17691 20591 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 22281 17731 22339 17737
rect 22281 17697 22293 17731
rect 22327 17728 22339 17731
rect 23474 17728 23480 17740
rect 22327 17700 23480 17728
rect 22327 17697 22339 17700
rect 22281 17691 22339 17697
rect 23474 17688 23480 17700
rect 23532 17688 23538 17740
rect 23842 17688 23848 17740
rect 23900 17688 23906 17740
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19352 17632 19901 17660
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 19889 17623 19947 17629
rect 22756 17632 23673 17660
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 13648 17564 13860 17592
rect 13648 17524 13676 17564
rect 11624 17496 13676 17524
rect 13832 17524 13860 17564
rect 13906 17552 13912 17604
rect 13964 17592 13970 17604
rect 15102 17592 15108 17604
rect 13964 17564 15108 17592
rect 13964 17552 13970 17564
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 15194 17552 15200 17604
rect 15252 17592 15258 17604
rect 15562 17592 15568 17604
rect 15252 17564 15568 17592
rect 15252 17552 15258 17564
rect 15562 17552 15568 17564
rect 15620 17552 15626 17604
rect 16500 17564 20024 17592
rect 16500 17524 16528 17564
rect 13832 17496 16528 17524
rect 17034 17484 17040 17536
rect 17092 17484 17098 17536
rect 17402 17484 17408 17536
rect 17460 17484 17466 17536
rect 17497 17527 17555 17533
rect 17497 17493 17509 17527
rect 17543 17524 17555 17527
rect 17862 17524 17868 17536
rect 17543 17496 17868 17524
rect 17543 17493 17555 17496
rect 17497 17487 17555 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19702 17524 19708 17536
rect 19475 17496 19708 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19794 17484 19800 17536
rect 19852 17484 19858 17536
rect 19996 17524 20024 17564
rect 20806 17552 20812 17604
rect 20864 17552 20870 17604
rect 20898 17552 20904 17604
rect 20956 17592 20962 17604
rect 20956 17564 21298 17592
rect 20956 17552 20962 17564
rect 22756 17536 22784 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 24578 17660 24584 17672
rect 23799 17632 24584 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 23382 17552 23388 17604
rect 23440 17592 23446 17604
rect 24765 17595 24823 17601
rect 24765 17592 24777 17595
rect 23440 17564 24777 17592
rect 23440 17552 23446 17564
rect 24765 17561 24777 17564
rect 24811 17561 24823 17595
rect 24765 17555 24823 17561
rect 22186 17524 22192 17536
rect 19996 17496 22192 17524
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 22738 17484 22744 17536
rect 22796 17484 22802 17536
rect 23293 17527 23351 17533
rect 23293 17493 23305 17527
rect 23339 17524 23351 17527
rect 24302 17524 24308 17536
rect 23339 17496 24308 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 24302 17484 24308 17496
rect 24360 17484 24366 17536
rect 24780 17524 24808 17555
rect 24946 17552 24952 17604
rect 25004 17552 25010 17604
rect 25409 17527 25467 17533
rect 25409 17524 25421 17527
rect 24780 17496 25421 17524
rect 25409 17493 25421 17496
rect 25455 17493 25467 17527
rect 25409 17487 25467 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6730 17320 6736 17332
rect 5951 17292 6736 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6730 17280 6736 17292
rect 6788 17280 6794 17332
rect 7193 17323 7251 17329
rect 7193 17289 7205 17323
rect 7239 17320 7251 17323
rect 8297 17323 8355 17329
rect 7239 17292 8248 17320
rect 7239 17289 7251 17292
rect 7193 17283 7251 17289
rect 5813 17255 5871 17261
rect 5813 17221 5825 17255
rect 5859 17252 5871 17255
rect 8220 17252 8248 17292
rect 8297 17289 8309 17323
rect 8343 17320 8355 17323
rect 8570 17320 8576 17332
rect 8343 17292 8576 17320
rect 8343 17289 8355 17292
rect 8297 17283 8355 17289
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 8662 17280 8668 17332
rect 8720 17280 8726 17332
rect 9766 17320 9772 17332
rect 9232 17292 9772 17320
rect 9232 17252 9260 17292
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10410 17320 10416 17332
rect 9916 17292 10416 17320
rect 9916 17280 9922 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 10560 17292 10903 17320
rect 10560 17280 10566 17292
rect 9674 17252 9680 17264
rect 5859 17224 7420 17252
rect 8220 17224 9260 17252
rect 9324 17224 9680 17252
rect 5859 17221 5871 17224
rect 5813 17215 5871 17221
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17184 3479 17187
rect 3970 17184 3976 17196
rect 3467 17156 3976 17184
rect 3467 17153 3479 17156
rect 3421 17147 3479 17153
rect 3970 17144 3976 17156
rect 4028 17184 4034 17196
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 4028 17156 4077 17184
rect 4028 17144 4034 17156
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 6086 17144 6092 17196
rect 6144 17144 6150 17196
rect 6362 17144 6368 17196
rect 6420 17184 6426 17196
rect 7392 17193 7420 17224
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6420 17156 6745 17184
rect 6420 17144 6426 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 7558 17184 7564 17196
rect 7423 17156 7564 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 7892 17156 8493 17184
rect 7892 17144 7898 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 8846 17144 8852 17196
rect 8904 17144 8910 17196
rect 9324 17193 9352 17224
rect 9674 17212 9680 17224
rect 9732 17212 9738 17264
rect 10875 17252 10903 17292
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 11020 17292 11069 17320
rect 11020 17280 11026 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 11057 17283 11115 17289
rect 12161 17323 12219 17329
rect 12161 17289 12173 17323
rect 12207 17320 12219 17323
rect 13817 17323 13875 17329
rect 12207 17292 13676 17320
rect 12207 17289 12219 17292
rect 12161 17283 12219 17289
rect 11146 17252 11152 17264
rect 10810 17224 11152 17252
rect 11146 17212 11152 17224
rect 11204 17252 11210 17264
rect 11204 17224 12388 17252
rect 11204 17212 11210 17224
rect 12360 17196 12388 17224
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11112 17156 12081 17184
rect 11112 17144 11118 17156
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12710 17184 12716 17196
rect 12400 17156 12716 17184
rect 12400 17144 12406 17156
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13648 17184 13676 17292
rect 13817 17289 13829 17323
rect 13863 17320 13875 17323
rect 17034 17320 17040 17332
rect 13863 17292 17040 17320
rect 13863 17289 13875 17292
rect 13817 17283 13875 17289
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 17218 17280 17224 17332
rect 17276 17280 17282 17332
rect 17313 17323 17371 17329
rect 17313 17289 17325 17323
rect 17359 17320 17371 17323
rect 17586 17320 17592 17332
rect 17359 17292 17592 17320
rect 17359 17289 17371 17292
rect 17313 17283 17371 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 20162 17320 20168 17332
rect 19392 17292 20168 17320
rect 19392 17280 19398 17292
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 22278 17320 22284 17332
rect 20864 17292 22284 17320
rect 20864 17280 20870 17292
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 23290 17320 23296 17332
rect 22428 17292 23296 17320
rect 22428 17280 22434 17292
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 23842 17280 23848 17332
rect 23900 17280 23906 17332
rect 13725 17255 13783 17261
rect 13725 17221 13737 17255
rect 13771 17252 13783 17255
rect 16666 17252 16672 17264
rect 13771 17224 16672 17252
rect 13771 17221 13783 17224
rect 13725 17215 13783 17221
rect 16666 17212 16672 17224
rect 16724 17212 16730 17264
rect 17402 17212 17408 17264
rect 17460 17252 17466 17264
rect 17770 17252 17776 17264
rect 17460 17224 17776 17252
rect 17460 17212 17466 17224
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 20346 17252 20352 17264
rect 19918 17224 20352 17252
rect 20180 17196 20208 17224
rect 20346 17212 20352 17224
rect 20404 17212 20410 17264
rect 20990 17212 20996 17264
rect 21048 17212 21054 17264
rect 25406 17252 25412 17264
rect 24228 17224 25412 17252
rect 14645 17187 14703 17193
rect 13648 17156 14044 17184
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 8205 17119 8263 17125
rect 6604 17088 8156 17116
rect 6604 17076 6610 17088
rect 3881 17051 3939 17057
rect 3881 17017 3893 17051
rect 3927 17048 3939 17051
rect 6822 17048 6828 17060
rect 3927 17020 6828 17048
rect 3927 17017 3939 17020
rect 3881 17011 3939 17017
rect 6822 17008 6828 17020
rect 6880 17008 6886 17060
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 4982 16980 4988 16992
rect 4939 16952 4988 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 6546 16940 6552 16992
rect 6604 16940 6610 16992
rect 8128 16980 8156 17088
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8864 17116 8892 17144
rect 8251 17088 8892 17116
rect 9585 17119 9643 17125
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 9585 17085 9597 17119
rect 9631 17116 9643 17119
rect 10870 17116 10876 17128
rect 9631 17088 10876 17116
rect 9631 17085 9643 17088
rect 9585 17079 9643 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 12032 17088 12265 17116
rect 12032 17076 12038 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 13906 17076 13912 17128
rect 13964 17076 13970 17128
rect 14016 17116 14044 17156
rect 14645 17153 14657 17187
rect 14691 17184 14703 17187
rect 14734 17184 14740 17196
rect 14691 17156 14740 17184
rect 14691 17153 14703 17156
rect 14645 17147 14703 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 15286 17144 15292 17196
rect 15344 17184 15350 17196
rect 15344 17156 15700 17184
rect 15344 17144 15350 17156
rect 15672 17116 15700 17156
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15896 17156 15945 17184
rect 15896 17144 15902 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 17862 17184 17868 17196
rect 15933 17147 15991 17153
rect 16040 17156 17868 17184
rect 16040 17125 16068 17156
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 20162 17144 20168 17196
rect 20220 17144 20226 17196
rect 20817 17191 20875 17197
rect 20817 17157 20829 17191
rect 20863 17188 20875 17191
rect 20863 17184 20944 17188
rect 21008 17184 21036 17212
rect 20863 17160 21036 17184
rect 20863 17157 20875 17160
rect 20817 17151 20875 17157
rect 20916 17156 21036 17160
rect 21450 17144 21456 17196
rect 21508 17144 21514 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 14016 17088 15608 17116
rect 15672 17088 16037 17116
rect 10594 17008 10600 17060
rect 10652 17048 10658 17060
rect 15580 17057 15608 17088
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16206 17076 16212 17128
rect 16264 17076 16270 17128
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17116 18751 17119
rect 20990 17116 20996 17128
rect 18739 17088 20996 17116
rect 18739 17085 18751 17088
rect 18693 17079 18751 17085
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 22020 17116 22048 17147
rect 22094 17144 22100 17196
rect 22152 17144 22158 17196
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 22373 17119 22431 17125
rect 22020 17088 22094 17116
rect 14829 17051 14887 17057
rect 14829 17048 14841 17051
rect 10652 17020 14841 17048
rect 10652 17008 10658 17020
rect 14829 17017 14841 17020
rect 14875 17017 14887 17051
rect 14829 17011 14887 17017
rect 15565 17051 15623 17057
rect 15565 17017 15577 17051
rect 15611 17017 15623 17051
rect 21910 17048 21916 17060
rect 15565 17011 15623 17017
rect 19720 17020 21916 17048
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 8128 16952 11713 16980
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 13354 16940 13360 16992
rect 13412 16940 13418 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16632 16952 16865 16980
rect 16632 16940 16638 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 19720 16980 19748 17020
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 17092 16952 19748 16980
rect 20625 16983 20683 16989
rect 17092 16940 17098 16952
rect 20625 16949 20637 16983
rect 20671 16980 20683 16983
rect 21174 16980 21180 16992
rect 20671 16952 21180 16980
rect 20671 16949 20683 16952
rect 20625 16943 20683 16949
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21726 16980 21732 16992
rect 21315 16952 21732 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 21818 16940 21824 16992
rect 21876 16940 21882 16992
rect 22066 16980 22094 17088
rect 22373 17085 22385 17119
rect 22419 17116 22431 17119
rect 24228 17116 24256 17224
rect 25406 17212 25412 17224
rect 25464 17212 25470 17264
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 22419 17088 24256 17116
rect 24320 17156 24961 17184
rect 22419 17085 22431 17088
rect 22373 17079 22431 17085
rect 23934 17048 23940 17060
rect 23400 17020 23940 17048
rect 23400 16980 23428 17020
rect 23934 17008 23940 17020
rect 23992 17008 23998 17060
rect 22066 16952 23428 16980
rect 23750 16940 23756 16992
rect 23808 16980 23814 16992
rect 24320 16989 24348 17156
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 25133 17051 25191 17057
rect 25133 17017 25145 17051
rect 25179 17048 25191 17051
rect 25406 17048 25412 17060
rect 25179 17020 25412 17048
rect 25179 17017 25191 17020
rect 25133 17011 25191 17017
rect 25406 17008 25412 17020
rect 25464 17008 25470 17060
rect 24305 16983 24363 16989
rect 24305 16980 24317 16983
rect 23808 16952 24317 16980
rect 23808 16940 23814 16952
rect 24305 16949 24317 16952
rect 24351 16949 24363 16983
rect 24305 16943 24363 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 4890 16736 4896 16788
rect 4948 16736 4954 16788
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 9950 16776 9956 16788
rect 5040 16748 9956 16776
rect 5040 16736 5046 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10689 16779 10747 16785
rect 10689 16776 10701 16779
rect 10284 16748 10701 16776
rect 10284 16736 10290 16748
rect 10689 16745 10701 16748
rect 10735 16745 10747 16779
rect 10689 16739 10747 16745
rect 11054 16736 11060 16788
rect 11112 16736 11118 16788
rect 11164 16748 15608 16776
rect 6730 16668 6736 16720
rect 6788 16668 6794 16720
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 9214 16708 9220 16720
rect 7524 16680 9220 16708
rect 7524 16668 7530 16680
rect 9214 16668 9220 16680
rect 9272 16668 9278 16720
rect 11164 16708 11192 16748
rect 10152 16680 11192 16708
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 6273 16575 6331 16581
rect 6273 16572 6285 16575
rect 5675 16544 6285 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 6273 16541 6285 16544
rect 6319 16572 6331 16575
rect 6748 16572 6776 16668
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16640 7435 16643
rect 7929 16643 7987 16649
rect 7423 16612 7880 16640
rect 7423 16609 7435 16612
rect 7377 16603 7435 16609
rect 6319 16544 6776 16572
rect 7852 16572 7880 16612
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 7975 16612 9628 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 7852 16544 8585 16572
rect 6319 16541 6331 16544
rect 6273 16535 6331 16541
rect 8573 16541 8585 16544
rect 8619 16572 8631 16575
rect 8938 16572 8944 16584
rect 8619 16544 8944 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 9600 16581 9628 16612
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 10152 16572 10180 16680
rect 14090 16668 14096 16720
rect 14148 16708 14154 16720
rect 15580 16708 15608 16748
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 19426 16776 19432 16788
rect 17644 16748 19432 16776
rect 17644 16736 17650 16748
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 19692 16779 19750 16785
rect 19692 16745 19704 16779
rect 19738 16776 19750 16779
rect 19738 16748 20760 16776
rect 19738 16745 19750 16748
rect 19692 16739 19750 16745
rect 17034 16708 17040 16720
rect 14148 16680 14412 16708
rect 15580 16680 17040 16708
rect 14148 16668 14154 16680
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11020 16612 11529 16640
rect 11020 16600 11026 16612
rect 11517 16609 11529 16612
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16640 12311 16643
rect 13722 16640 13728 16652
rect 12299 16612 13728 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14274 16600 14280 16652
rect 14332 16600 14338 16652
rect 14384 16640 14412 16680
rect 17034 16668 17040 16680
rect 17092 16668 17098 16720
rect 20732 16708 20760 16748
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 21048 16748 21189 16776
rect 21048 16736 21054 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 21177 16739 21235 16745
rect 21358 16708 21364 16720
rect 20732 16680 21364 16708
rect 21358 16668 21364 16680
rect 21416 16668 21422 16720
rect 14550 16640 14556 16652
rect 14384 16612 14556 16640
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 16850 16600 16856 16652
rect 16908 16640 16914 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 16908 16612 17141 16640
rect 16908 16600 16914 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 19334 16640 19340 16652
rect 17451 16612 19340 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 22094 16640 22100 16652
rect 19475 16612 22100 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 22094 16600 22100 16612
rect 22152 16640 22158 16652
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 22152 16612 22293 16640
rect 22152 16600 22158 16612
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 22281 16603 22339 16609
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 23566 16640 23572 16652
rect 22603 16612 23572 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 24857 16643 24915 16649
rect 24857 16640 24869 16643
rect 24636 16612 24869 16640
rect 24636 16600 24642 16612
rect 24857 16609 24869 16612
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 9631 16544 10180 16572
rect 10229 16575 10287 16581
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 10229 16541 10241 16575
rect 10275 16572 10287 16575
rect 11054 16572 11060 16584
rect 10275 16544 11060 16572
rect 10275 16541 10287 16544
rect 10229 16535 10287 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 21818 16532 21824 16584
rect 21876 16532 21882 16584
rect 5166 16464 5172 16516
rect 5224 16504 5230 16516
rect 12526 16504 12532 16516
rect 5224 16476 12532 16504
rect 5224 16464 5230 16476
rect 12526 16464 12532 16476
rect 12584 16464 12590 16516
rect 12710 16464 12716 16516
rect 12768 16464 12774 16516
rect 15286 16464 15292 16516
rect 15344 16464 15350 16516
rect 17862 16464 17868 16516
rect 17920 16464 17926 16516
rect 18690 16464 18696 16516
rect 18748 16504 18754 16516
rect 20162 16504 20168 16516
rect 18748 16476 20168 16504
rect 18748 16464 18754 16476
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 23566 16464 23572 16516
rect 23624 16464 23630 16516
rect 24670 16464 24676 16516
rect 24728 16464 24734 16516
rect 6086 16396 6092 16448
rect 6144 16396 6150 16448
rect 8386 16396 8392 16448
rect 8444 16396 8450 16448
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9950 16436 9956 16448
rect 9447 16408 9956 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10042 16396 10048 16448
rect 10100 16396 10106 16448
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12124 16408 13737 16436
rect 12124 16396 12130 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 17310 16396 17316 16448
rect 17368 16436 17374 16448
rect 18877 16439 18935 16445
rect 18877 16436 18889 16439
rect 17368 16408 18889 16436
rect 17368 16396 17374 16408
rect 18877 16405 18889 16408
rect 18923 16436 18935 16439
rect 21266 16436 21272 16448
rect 18923 16408 21272 16436
rect 18923 16405 18935 16408
rect 18877 16399 18935 16405
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 21450 16396 21456 16448
rect 21508 16436 21514 16448
rect 22002 16436 22008 16448
rect 21508 16408 22008 16436
rect 21508 16396 21514 16408
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 23934 16396 23940 16448
rect 23992 16436 23998 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23992 16408 24041 16436
rect 23992 16396 23998 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 9122 16192 9128 16244
rect 9180 16192 9186 16244
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 9272 16204 10609 16232
rect 9272 16192 9278 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 10962 16192 10968 16244
rect 11020 16192 11026 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 11572 16204 13461 16232
rect 11572 16192 11578 16204
rect 13449 16201 13461 16204
rect 13495 16232 13507 16235
rect 16206 16232 16212 16244
rect 13495 16204 16212 16232
rect 13495 16201 13507 16204
rect 13449 16195 13507 16201
rect 16206 16192 16212 16204
rect 16264 16192 16270 16244
rect 18506 16192 18512 16244
rect 18564 16192 18570 16244
rect 18966 16192 18972 16244
rect 19024 16232 19030 16244
rect 19242 16232 19248 16244
rect 19024 16204 19248 16232
rect 19024 16192 19030 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19429 16235 19487 16241
rect 19429 16201 19441 16235
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 11054 16164 11060 16176
rect 9876 16136 11060 16164
rect 5166 16056 5172 16108
rect 5224 16056 5230 16108
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 8570 16096 8576 16108
rect 8527 16068 8576 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 4246 15988 4252 16040
rect 4304 16028 4310 16040
rect 5445 16031 5503 16037
rect 5445 16028 5457 16031
rect 4304 16000 5457 16028
rect 4304 15988 4310 16000
rect 5445 15997 5457 16000
rect 5491 15997 5503 16031
rect 5445 15991 5503 15997
rect 9033 16031 9091 16037
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9876 16028 9904 16136
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 11977 16167 12035 16173
rect 11977 16133 11989 16167
rect 12023 16164 12035 16167
rect 12066 16164 12072 16176
rect 12023 16136 12072 16164
rect 12023 16133 12035 16136
rect 11977 16127 12035 16133
rect 12066 16124 12072 16136
rect 12124 16124 12130 16176
rect 12250 16124 12256 16176
rect 12308 16164 12314 16176
rect 12434 16164 12440 16176
rect 12308 16136 12440 16164
rect 12308 16124 12314 16136
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 14369 16167 14427 16173
rect 14369 16133 14381 16167
rect 14415 16164 14427 16167
rect 19444 16164 19472 16195
rect 19886 16192 19892 16244
rect 19944 16192 19950 16244
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16232 21143 16235
rect 21818 16232 21824 16244
rect 21131 16204 21824 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 22002 16192 22008 16244
rect 22060 16232 22066 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 22060 16204 22477 16232
rect 22060 16192 22066 16204
rect 22465 16201 22477 16204
rect 22511 16201 22523 16235
rect 22465 16195 22523 16201
rect 23845 16235 23903 16241
rect 23845 16201 23857 16235
rect 23891 16232 23903 16235
rect 24394 16232 24400 16244
rect 23891 16204 24400 16232
rect 23891 16201 23903 16204
rect 23845 16195 23903 16201
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 14415 16136 19472 16164
rect 14415 16133 14427 16136
rect 14369 16127 14427 16133
rect 20438 16124 20444 16176
rect 20496 16164 20502 16176
rect 21177 16167 21235 16173
rect 21177 16164 21189 16167
rect 20496 16136 21189 16164
rect 20496 16124 20502 16136
rect 21177 16133 21189 16136
rect 21223 16133 21235 16167
rect 21177 16127 21235 16133
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 10226 16096 10232 16108
rect 9999 16068 10232 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 14090 16056 14096 16108
rect 14148 16096 14154 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 14148 16068 14289 16096
rect 14148 16056 14154 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15896 16068 15945 16096
rect 15896 16056 15902 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 17126 16056 17132 16108
rect 17184 16096 17190 16108
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 17184 16068 17233 16096
rect 17184 16056 17190 16068
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18690 16096 18696 16108
rect 18012 16068 18696 16096
rect 18012 16056 18018 16068
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 9079 16000 9904 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 10192 16000 10425 16028
rect 10192 15988 10198 16000
rect 10413 15997 10425 16000
rect 10459 16028 10471 16031
rect 10502 16028 10508 16040
rect 10459 16000 10508 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 10652 16000 10916 16028
rect 10652 15988 10658 16000
rect 6086 15920 6092 15972
rect 6144 15960 6150 15972
rect 10888 15960 10916 16000
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 11020 16000 11069 16028
rect 11020 15988 11026 16000
rect 11057 15997 11069 16000
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 12066 16028 12072 16040
rect 11808 16000 12072 16028
rect 11808 15960 11836 16000
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 16025 16031 16083 16037
rect 16025 16028 16037 16031
rect 15712 16000 16037 16028
rect 15712 15988 15718 16000
rect 16025 15997 16037 16000
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 15997 16175 16031
rect 16117 15991 16175 15997
rect 6144 15932 10732 15960
rect 10888 15932 11836 15960
rect 6144 15920 6150 15932
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 10594 15892 10600 15904
rect 7064 15864 10600 15892
rect 7064 15852 7070 15864
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 10704 15892 10732 15932
rect 15562 15920 15568 15972
rect 15620 15920 15626 15972
rect 13814 15892 13820 15904
rect 10704 15864 13820 15892
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 16132 15892 16160 15991
rect 16758 15988 16764 16040
rect 16816 16028 16822 16040
rect 19812 16028 19840 16059
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 21048 16068 21312 16096
rect 21048 16056 21054 16068
rect 16816 16000 19840 16028
rect 16816 15988 16822 16000
rect 20070 15988 20076 16040
rect 20128 15988 20134 16040
rect 21284 16037 21312 16068
rect 21634 16056 21640 16108
rect 21692 16096 21698 16108
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 21692 16068 22385 16096
rect 21692 16056 21698 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16096 23811 16099
rect 24210 16096 24216 16108
rect 23799 16068 24216 16096
rect 23799 16065 23811 16068
rect 23753 16059 23811 16065
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 24670 16056 24676 16108
rect 24728 16056 24734 16108
rect 21269 16031 21327 16037
rect 21269 15997 21281 16031
rect 21315 15997 21327 16031
rect 21269 15991 21327 15997
rect 22278 15988 22284 16040
rect 22336 16028 22342 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22336 16000 22569 16028
rect 22336 15988 22342 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 23934 15988 23940 16040
rect 23992 15988 23998 16040
rect 17034 15920 17040 15972
rect 17092 15960 17098 15972
rect 24857 15963 24915 15969
rect 17092 15932 24808 15960
rect 17092 15920 17098 15932
rect 14700 15864 16160 15892
rect 14700 15852 14706 15864
rect 18966 15852 18972 15904
rect 19024 15892 19030 15904
rect 20717 15895 20775 15901
rect 20717 15892 20729 15895
rect 19024 15864 20729 15892
rect 19024 15852 19030 15864
rect 20717 15861 20729 15864
rect 20763 15861 20775 15895
rect 20717 15855 20775 15861
rect 21634 15852 21640 15904
rect 21692 15892 21698 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21692 15864 22017 15892
rect 21692 15852 21698 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 22370 15852 22376 15904
rect 22428 15892 22434 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 22428 15864 23397 15892
rect 22428 15852 22434 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 24780 15892 24808 15932
rect 24857 15929 24869 15963
rect 24903 15960 24915 15963
rect 25222 15960 25228 15972
rect 24903 15932 25228 15960
rect 24903 15929 24915 15932
rect 24857 15923 24915 15929
rect 25222 15920 25228 15932
rect 25280 15920 25286 15972
rect 25130 15892 25136 15904
rect 24780 15864 25136 15892
rect 23385 15855 23443 15861
rect 25130 15852 25136 15864
rect 25188 15852 25194 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 13906 15688 13912 15700
rect 8536 15660 13912 15688
rect 8536 15648 8542 15660
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 16025 15691 16083 15697
rect 16025 15688 16037 15691
rect 15160 15660 16037 15688
rect 15160 15648 15166 15660
rect 16025 15657 16037 15660
rect 16071 15657 16083 15691
rect 16025 15651 16083 15657
rect 18782 15648 18788 15700
rect 18840 15648 18846 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 22462 15688 22468 15700
rect 20763 15660 22468 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 9493 15623 9551 15629
rect 9493 15589 9505 15623
rect 9539 15620 9551 15623
rect 10226 15620 10232 15632
rect 9539 15592 10232 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 12713 15623 12771 15629
rect 12713 15620 12725 15623
rect 12124 15592 12725 15620
rect 12124 15580 12130 15592
rect 12713 15589 12725 15592
rect 12759 15589 12771 15623
rect 12713 15583 12771 15589
rect 19521 15623 19579 15629
rect 19521 15589 19533 15623
rect 19567 15620 19579 15623
rect 19978 15620 19984 15632
rect 19567 15592 19984 15620
rect 19567 15589 19579 15592
rect 19521 15583 19579 15589
rect 19978 15580 19984 15592
rect 20036 15580 20042 15632
rect 22554 15620 22560 15632
rect 21192 15592 22560 15620
rect 9401 15555 9459 15561
rect 9401 15521 9413 15555
rect 9447 15552 9459 15555
rect 10965 15555 11023 15561
rect 9447 15524 10548 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 10520 15496 10548 15524
rect 10965 15521 10977 15555
rect 11011 15552 11023 15555
rect 11514 15552 11520 15564
rect 11011 15524 11520 15552
rect 11011 15521 11023 15524
rect 10965 15515 11023 15521
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 13722 15552 13728 15564
rect 13403 15524 13728 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15552 14611 15555
rect 16482 15552 16488 15564
rect 14599 15524 16488 15552
rect 14599 15521 14611 15524
rect 14553 15515 14611 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 17310 15512 17316 15564
rect 17368 15512 17374 15564
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15552 20223 15555
rect 20254 15552 20260 15564
rect 20211 15524 20260 15552
rect 20211 15521 20223 15524
rect 20165 15515 20223 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 21192 15561 21220 15592
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 21177 15555 21235 15561
rect 21177 15521 21189 15555
rect 21223 15521 21235 15555
rect 21177 15515 21235 15521
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 24765 15555 24823 15561
rect 24765 15552 24777 15555
rect 22066 15524 24777 15552
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15484 9735 15487
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9723 15456 10241 15484
rect 9723 15453 9735 15456
rect 9677 15447 9735 15453
rect 10229 15453 10241 15456
rect 10275 15484 10287 15487
rect 10318 15484 10324 15496
rect 10275 15456 10324 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 10686 15444 10692 15496
rect 10744 15444 10750 15496
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20530 15484 20536 15496
rect 19935 15456 20536 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 22066 15484 22094 15524
rect 24765 15521 24777 15524
rect 24811 15521 24823 15555
rect 24765 15515 24823 15521
rect 21131 15456 22094 15484
rect 22189 15487 22247 15493
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 22189 15453 22201 15487
rect 22235 15484 22247 15487
rect 22278 15484 22284 15496
rect 22235 15456 22284 15484
rect 22235 15453 22247 15456
rect 22189 15447 22247 15453
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 23658 15484 23664 15496
rect 23615 15456 23664 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 12342 15416 12348 15428
rect 12190 15388 12348 15416
rect 12342 15376 12348 15388
rect 12400 15376 12406 15428
rect 13081 15419 13139 15425
rect 13081 15385 13093 15419
rect 13127 15416 13139 15419
rect 13354 15416 13360 15428
rect 13127 15388 13360 15416
rect 13127 15385 13139 15388
rect 13081 15379 13139 15385
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 15286 15376 15292 15428
rect 15344 15376 15350 15428
rect 17310 15376 17316 15428
rect 17368 15416 17374 15428
rect 17770 15416 17776 15428
rect 17368 15388 17776 15416
rect 17368 15376 17374 15388
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 19794 15376 19800 15428
rect 19852 15416 19858 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19852 15388 19993 15416
rect 19852 15376 19858 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 21174 15376 21180 15428
rect 21232 15416 21238 15428
rect 22005 15419 22063 15425
rect 22005 15416 22017 15419
rect 21232 15388 22017 15416
rect 21232 15376 21238 15388
rect 22005 15385 22017 15388
rect 22051 15385 22063 15419
rect 22005 15379 22063 15385
rect 22741 15419 22799 15425
rect 22741 15385 22753 15419
rect 22787 15385 22799 15419
rect 22741 15379 22799 15385
rect 10321 15351 10379 15357
rect 10321 15317 10333 15351
rect 10367 15348 10379 15351
rect 11790 15348 11796 15360
rect 10367 15320 11796 15348
rect 10367 15317 10379 15320
rect 10321 15311 10379 15317
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12437 15351 12495 15357
rect 12437 15348 12449 15351
rect 12032 15320 12449 15348
rect 12032 15308 12038 15320
rect 12437 15317 12449 15320
rect 12483 15317 12495 15351
rect 12437 15311 12495 15317
rect 13173 15351 13231 15357
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 16574 15348 16580 15360
rect 13219 15320 16580 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 19886 15348 19892 15360
rect 17276 15320 19892 15348
rect 17276 15308 17282 15320
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 21726 15308 21732 15360
rect 21784 15348 21790 15360
rect 22756 15348 22784 15379
rect 21784 15320 22784 15348
rect 21784 15308 21790 15320
rect 22830 15308 22836 15360
rect 22888 15308 22894 15360
rect 23290 15308 23296 15360
rect 23348 15348 23354 15360
rect 23385 15351 23443 15357
rect 23385 15348 23397 15351
rect 23348 15320 23397 15348
rect 23348 15308 23354 15320
rect 23385 15317 23397 15320
rect 23431 15317 23443 15351
rect 23385 15311 23443 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 12066 15144 12072 15156
rect 11296 15116 12072 15144
rect 11296 15104 11302 15116
rect 12066 15104 12072 15116
rect 12124 15144 12130 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12124 15116 13461 15144
rect 12124 15104 12130 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 14829 15147 14887 15153
rect 14829 15113 14841 15147
rect 14875 15144 14887 15147
rect 15378 15144 15384 15156
rect 14875 15116 15384 15144
rect 14875 15113 14887 15116
rect 14829 15107 14887 15113
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 16758 15144 16764 15156
rect 15519 15116 16764 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 16850 15104 16856 15156
rect 16908 15144 16914 15156
rect 21177 15147 21235 15153
rect 16908 15116 19472 15144
rect 16908 15104 16914 15116
rect 10505 15079 10563 15085
rect 10505 15045 10517 15079
rect 10551 15076 10563 15079
rect 11882 15076 11888 15088
rect 10551 15048 11888 15076
rect 10551 15045 10563 15048
rect 10505 15039 10563 15045
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 10778 15008 10784 15020
rect 9907 14980 10784 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 11164 15017 11192 15048
rect 11882 15036 11888 15048
rect 11940 15036 11946 15088
rect 12434 15036 12440 15088
rect 12492 15036 12498 15088
rect 13906 15036 13912 15088
rect 13964 15076 13970 15088
rect 17218 15076 17224 15088
rect 13964 15048 17224 15076
rect 13964 15036 13970 15048
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 17770 15036 17776 15088
rect 17828 15036 17834 15088
rect 19444 15020 19472 15116
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 21358 15144 21364 15156
rect 21223 15116 21364 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 24670 15104 24676 15156
rect 24728 15144 24734 15156
rect 25038 15144 25044 15156
rect 24728 15116 25044 15144
rect 24728 15104 24734 15116
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 25130 15104 25136 15156
rect 25188 15104 25194 15156
rect 20990 15076 20996 15088
rect 20930 15048 20996 15076
rect 20990 15036 20996 15048
rect 21048 15076 21054 15088
rect 21266 15076 21272 15088
rect 21048 15048 21272 15076
rect 21048 15036 21054 15048
rect 21266 15036 21272 15048
rect 21324 15036 21330 15088
rect 22097 15079 22155 15085
rect 22097 15045 22109 15079
rect 22143 15076 22155 15079
rect 22646 15076 22652 15088
rect 22143 15048 22652 15076
rect 22143 15045 22155 15048
rect 22097 15039 22155 15045
rect 22646 15036 22652 15048
rect 22704 15036 22710 15088
rect 23658 15036 23664 15088
rect 23716 15036 23722 15088
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15059 14980 15424 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11698 14940 11704 14952
rect 10744 14912 11704 14940
rect 10744 14900 10750 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12434 14940 12440 14952
rect 12023 14912 12440 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12434 14900 12440 14912
rect 12492 14940 12498 14952
rect 14642 14940 14648 14952
rect 12492 14912 14648 14940
rect 12492 14900 12498 14912
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 15396 14872 15424 14980
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 15764 14980 16313 15008
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 15764 14940 15792 14980
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 19426 14968 19432 15020
rect 19484 14968 19490 15020
rect 25314 14968 25320 15020
rect 25372 14968 25378 15020
rect 15528 14912 15792 14940
rect 17129 14943 17187 14949
rect 15528 14900 15534 14912
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 18782 14940 18788 14952
rect 17175 14912 18788 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 19702 14900 19708 14952
rect 19760 14900 19766 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22925 14943 22983 14949
rect 22925 14940 22937 14943
rect 21968 14912 22937 14940
rect 21968 14900 21974 14912
rect 22925 14909 22937 14912
rect 22971 14909 22983 14943
rect 22925 14903 22983 14909
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14940 23259 14943
rect 23934 14940 23940 14952
rect 23247 14912 23940 14940
rect 23247 14909 23259 14912
rect 23201 14903 23259 14909
rect 23934 14900 23940 14912
rect 23992 14900 23998 14952
rect 16666 14872 16672 14884
rect 15396 14844 16672 14872
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 18874 14872 18880 14884
rect 18524 14844 18880 14872
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 16117 14807 16175 14813
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 18524 14804 18552 14844
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 22281 14875 22339 14881
rect 22281 14841 22293 14875
rect 22327 14872 22339 14875
rect 22462 14872 22468 14884
rect 22327 14844 22468 14872
rect 22327 14841 22339 14844
rect 22281 14835 22339 14841
rect 22462 14832 22468 14844
rect 22520 14832 22526 14884
rect 16163 14776 18552 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 10652 14572 12020 14600
rect 10652 14560 10658 14572
rect 11992 14532 12020 14572
rect 12434 14560 12440 14612
rect 12492 14560 12498 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 12860 14572 12909 14600
rect 12860 14560 12866 14572
rect 12897 14569 12909 14572
rect 12943 14569 12955 14603
rect 12897 14563 12955 14569
rect 13265 14603 13323 14609
rect 13265 14569 13277 14603
rect 13311 14600 13323 14603
rect 13354 14600 13360 14612
rect 13311 14572 13360 14600
rect 13311 14569 13323 14572
rect 13265 14563 13323 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 15010 14600 15016 14612
rect 13872 14572 15016 14600
rect 13872 14560 13878 14572
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 23382 14600 23388 14612
rect 15712 14572 23388 14600
rect 15712 14560 15718 14572
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 13998 14532 14004 14544
rect 11992 14504 14004 14532
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 16025 14535 16083 14541
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 16482 14532 16488 14544
rect 16071 14504 16488 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 16482 14492 16488 14504
rect 16540 14492 16546 14544
rect 18233 14535 18291 14541
rect 18233 14501 18245 14535
rect 18279 14532 18291 14535
rect 18322 14532 18328 14544
rect 18279 14504 18328 14532
rect 18279 14501 18291 14504
rect 18233 14495 18291 14501
rect 18322 14492 18328 14504
rect 18380 14532 18386 14544
rect 18782 14532 18788 14544
rect 18380 14504 18788 14532
rect 18380 14492 18386 14504
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14532 19487 14535
rect 21174 14532 21180 14544
rect 19475 14504 21180 14532
rect 19475 14501 19487 14504
rect 19429 14495 19487 14501
rect 21174 14492 21180 14504
rect 21232 14492 21238 14544
rect 23293 14535 23351 14541
rect 23293 14532 23305 14535
rect 22066 14504 23305 14532
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11974 14464 11980 14476
rect 11011 14436 11980 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 16761 14467 16819 14473
rect 14332 14436 16528 14464
rect 14332 14424 14338 14436
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 16500 14405 16528 14436
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 18598 14464 18604 14476
rect 16807 14436 18604 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 18598 14424 18604 14436
rect 18656 14464 18662 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 18656 14436 19993 14464
rect 18656 14424 18662 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 18923 14368 19809 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 12342 14328 12348 14340
rect 12190 14300 12348 14328
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 14550 14288 14556 14340
rect 14608 14288 14614 14340
rect 15286 14288 15292 14340
rect 15344 14288 15350 14340
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 14826 14260 14832 14272
rect 12768 14232 14832 14260
rect 12768 14220 12774 14232
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 16500 14260 16528 14359
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 22066 14396 22094 14504
rect 23293 14501 23305 14504
rect 23339 14501 23351 14535
rect 23293 14495 23351 14501
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24026 14464 24032 14476
rect 23983 14436 24032 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24026 14424 24032 14436
rect 24084 14424 24090 14476
rect 19944 14368 22094 14396
rect 23661 14399 23719 14405
rect 19944 14356 19950 14368
rect 23661 14365 23673 14399
rect 23707 14396 23719 14399
rect 25038 14396 25044 14408
rect 23707 14368 25044 14396
rect 23707 14365 23719 14368
rect 23661 14359 23719 14365
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 16724 14300 17172 14328
rect 16724 14288 16730 14300
rect 17034 14260 17040 14272
rect 16500 14232 17040 14260
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 17144 14260 17172 14300
rect 17310 14288 17316 14340
rect 17368 14288 17374 14340
rect 18506 14288 18512 14340
rect 18564 14328 18570 14340
rect 20809 14331 20867 14337
rect 20809 14328 20821 14331
rect 18564 14300 20821 14328
rect 18564 14288 18570 14300
rect 20809 14297 20821 14300
rect 20855 14297 20867 14331
rect 20809 14291 20867 14297
rect 20898 14288 20904 14340
rect 20956 14328 20962 14340
rect 23566 14328 23572 14340
rect 20956 14300 23572 14328
rect 20956 14288 20962 14300
rect 23566 14288 23572 14300
rect 23624 14288 23630 14340
rect 23753 14331 23811 14337
rect 23753 14297 23765 14331
rect 23799 14328 23811 14331
rect 24486 14328 24492 14340
rect 23799 14300 24492 14328
rect 23799 14297 23811 14300
rect 23753 14291 23811 14297
rect 24486 14288 24492 14300
rect 24544 14288 24550 14340
rect 24673 14331 24731 14337
rect 24673 14297 24685 14331
rect 24719 14328 24731 14331
rect 25590 14328 25596 14340
rect 24719 14300 25596 14328
rect 24719 14297 24731 14300
rect 24673 14291 24731 14297
rect 25590 14288 25596 14300
rect 25648 14288 25654 14340
rect 19058 14260 19064 14272
rect 17144 14232 19064 14260
rect 19058 14220 19064 14232
rect 19116 14220 19122 14272
rect 19518 14220 19524 14272
rect 19576 14260 19582 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19576 14232 19901 14260
rect 19576 14220 19582 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 21910 14220 21916 14272
rect 21968 14260 21974 14272
rect 22097 14263 22155 14269
rect 22097 14260 22109 14263
rect 21968 14232 22109 14260
rect 21968 14220 21974 14232
rect 22097 14229 22109 14232
rect 22143 14229 22155 14263
rect 22097 14223 22155 14229
rect 23842 14220 23848 14272
rect 23900 14260 23906 14272
rect 24765 14263 24823 14269
rect 24765 14260 24777 14263
rect 23900 14232 24777 14260
rect 23900 14220 23906 14232
rect 24765 14229 24777 14232
rect 24811 14229 24823 14263
rect 24765 14223 24823 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13446 14056 13452 14068
rect 13219 14028 13452 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 14182 14056 14188 14068
rect 13556 14028 14188 14056
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 13556 13988 13584 14028
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 14608 14028 15761 14056
rect 14608 14016 14614 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 15896 14028 16129 14056
rect 15896 14016 15902 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17218 14056 17224 14068
rect 17083 14028 17224 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 17678 14056 17684 14068
rect 17543 14028 17684 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19484 14028 19533 14056
rect 19484 14016 19490 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20717 14059 20775 14065
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 20990 14056 20996 14068
rect 20763 14028 20996 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21085 14059 21143 14065
rect 21085 14025 21097 14059
rect 21131 14056 21143 14059
rect 23474 14056 23480 14068
rect 21131 14028 23480 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 23566 14016 23572 14068
rect 23624 14056 23630 14068
rect 25225 14059 25283 14065
rect 25225 14056 25237 14059
rect 23624 14028 25237 14056
rect 23624 14016 23630 14028
rect 25225 14025 25237 14028
rect 25271 14025 25283 14059
rect 25225 14019 25283 14025
rect 12299 13960 13584 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 12802 13920 12808 13932
rect 12575 13892 12808 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 12912 13929 12940 13960
rect 13814 13948 13820 14000
rect 13872 13948 13878 14000
rect 14274 13988 14280 14000
rect 14016 13960 14280 13988
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13832 13920 13860 13948
rect 14016 13929 14044 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 15286 13948 15292 14000
rect 15344 13948 15350 14000
rect 17586 13988 17592 14000
rect 16316 13960 17592 13988
rect 16316 13929 16344 13960
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 18233 13991 18291 13997
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18322 13988 18328 14000
rect 18279 13960 18328 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18322 13948 18328 13960
rect 18380 13988 18386 14000
rect 18506 13988 18512 14000
rect 18380 13960 18512 13988
rect 18380 13948 18386 13960
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 20898 13988 20904 14000
rect 19116 13960 20904 13988
rect 19116 13948 19122 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21177 13991 21235 13997
rect 21177 13988 21189 13991
rect 21008 13960 21189 13988
rect 13403 13892 13860 13920
rect 14001 13923 14059 13929
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 14001 13889 14013 13923
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 16482 13880 16488 13932
rect 16540 13920 16546 13932
rect 17310 13920 17316 13932
rect 16540 13892 17316 13920
rect 16540 13880 16546 13892
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 18414 13920 18420 13932
rect 17451 13892 18420 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21008 13920 21036 13960
rect 21177 13957 21189 13960
rect 21223 13957 21235 13991
rect 21177 13951 21235 13957
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 20772 13892 21036 13920
rect 21100 13892 22017 13920
rect 20772 13880 20778 13892
rect 13906 13852 13912 13864
rect 12360 13824 13912 13852
rect 12360 13793 12388 13824
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 17586 13852 17592 13864
rect 14424 13824 17592 13852
rect 14424 13812 14430 13824
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 12345 13787 12403 13793
rect 12345 13753 12357 13787
rect 12391 13753 12403 13787
rect 12345 13747 12403 13753
rect 16022 13744 16028 13796
rect 16080 13784 16086 13796
rect 17696 13784 17724 13815
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 21100 13852 21128 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 23658 13880 23664 13932
rect 23716 13880 23722 13932
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 17828 13824 21128 13852
rect 21269 13855 21327 13861
rect 17828 13812 17834 13824
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 21269 13815 21327 13821
rect 16080 13756 17724 13784
rect 16080 13744 16086 13756
rect 14264 13719 14322 13725
rect 14264 13685 14276 13719
rect 14310 13716 14322 13719
rect 15562 13716 15568 13728
rect 14310 13688 15568 13716
rect 14310 13685 14322 13688
rect 14264 13679 14322 13685
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 17696 13716 17724 13756
rect 19702 13744 19708 13796
rect 19760 13784 19766 13796
rect 21284 13784 21312 13815
rect 21910 13812 21916 13864
rect 21968 13852 21974 13864
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 21968 13824 22293 13852
rect 21968 13812 21974 13824
rect 22281 13821 22293 13824
rect 22327 13821 22339 13855
rect 22281 13815 22339 13821
rect 24026 13812 24032 13864
rect 24084 13812 24090 13864
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 25148 13852 25176 13883
rect 24544 13824 25176 13852
rect 24544 13812 24550 13824
rect 21450 13784 21456 13796
rect 19760 13756 21456 13784
rect 19760 13744 19766 13756
rect 21450 13744 21456 13756
rect 21508 13744 21514 13796
rect 21542 13744 21548 13796
rect 21600 13784 21606 13796
rect 22186 13784 22192 13796
rect 21600 13756 22192 13784
rect 21600 13744 21606 13756
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 20162 13716 20168 13728
rect 17696 13688 20168 13716
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 21358 13716 21364 13728
rect 20404 13688 21364 13716
rect 20404 13676 20410 13688
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 21726 13676 21732 13728
rect 21784 13716 21790 13728
rect 22097 13719 22155 13725
rect 22097 13716 22109 13719
rect 21784 13688 22109 13716
rect 21784 13676 21790 13688
rect 22097 13685 22109 13688
rect 22143 13685 22155 13719
rect 22097 13679 22155 13685
rect 22544 13719 22602 13725
rect 22544 13685 22556 13719
rect 22590 13716 22602 13719
rect 24670 13716 24676 13728
rect 22590 13688 24676 13716
rect 22590 13685 22602 13688
rect 22544 13679 22602 13685
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13228 13484 13553 13512
rect 13228 13472 13234 13484
rect 13541 13481 13553 13484
rect 13587 13512 13599 13515
rect 17402 13512 17408 13524
rect 13587 13484 17408 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 18233 13515 18291 13521
rect 18233 13481 18245 13515
rect 18279 13512 18291 13515
rect 18874 13512 18880 13524
rect 18279 13484 18880 13512
rect 18279 13481 18291 13484
rect 18233 13475 18291 13481
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 20070 13512 20076 13524
rect 18984 13484 20076 13512
rect 15562 13404 15568 13456
rect 15620 13444 15626 13456
rect 16025 13447 16083 13453
rect 16025 13444 16037 13447
rect 15620 13416 16037 13444
rect 15620 13404 15626 13416
rect 16025 13413 16037 13416
rect 16071 13444 16083 13447
rect 18984 13444 19012 13484
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 21450 13472 21456 13524
rect 21508 13472 21514 13524
rect 16071 13416 19012 13444
rect 24581 13447 24639 13453
rect 16071 13413 16083 13416
rect 16025 13407 16083 13413
rect 24581 13413 24593 13447
rect 24627 13413 24639 13447
rect 24581 13407 24639 13413
rect 12066 13336 12072 13388
rect 12124 13336 12130 13388
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 19150 13376 19156 13388
rect 17000 13348 19156 13376
rect 17000 13336 17006 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19484 13348 19717 13376
rect 19484 13336 19490 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13376 20039 13379
rect 20346 13376 20352 13388
rect 20027 13348 20352 13376
rect 20027 13345 20039 13348
rect 19981 13339 20039 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 24596 13376 24624 13407
rect 20588 13348 24624 13376
rect 20588 13336 20594 13348
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 25041 13379 25099 13385
rect 25041 13376 25053 13379
rect 24912 13348 25053 13376
rect 24912 13336 24918 13348
rect 25041 13345 25053 13348
rect 25087 13345 25099 13379
rect 25041 13339 25099 13345
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 9582 13268 9588 13320
rect 9640 13268 9646 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 10888 13280 11805 13308
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10686 13172 10692 13184
rect 10192 13144 10692 13172
rect 10192 13132 10198 13144
rect 10686 13132 10692 13144
rect 10744 13172 10750 13184
rect 10888 13181 10916 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 21910 13268 21916 13320
rect 21968 13268 21974 13320
rect 12452 13212 12558 13240
rect 12452 13184 12480 13212
rect 13722 13200 13728 13252
rect 13780 13240 13786 13252
rect 14553 13243 14611 13249
rect 14553 13240 14565 13243
rect 13780 13212 14565 13240
rect 13780 13200 13786 13212
rect 14553 13209 14565 13212
rect 14599 13240 14611 13243
rect 14642 13240 14648 13252
rect 14599 13212 14648 13240
rect 14599 13209 14611 13212
rect 14553 13203 14611 13209
rect 14642 13200 14648 13212
rect 14700 13200 14706 13252
rect 16482 13240 16488 13252
rect 14936 13212 15042 13240
rect 16224 13212 16488 13240
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 13630 13172 13636 13184
rect 12492 13144 13636 13172
rect 12492 13132 12498 13144
rect 13630 13132 13636 13144
rect 13688 13172 13694 13184
rect 14936 13172 14964 13212
rect 15286 13172 15292 13184
rect 13688 13144 15292 13172
rect 13688 13132 13694 13144
rect 15286 13132 15292 13144
rect 15344 13172 15350 13184
rect 16224 13172 16252 13212
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 19150 13240 19156 13252
rect 19024 13212 19156 13240
rect 19024 13200 19030 13212
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 21266 13240 21272 13252
rect 21206 13212 21272 13240
rect 21266 13200 21272 13212
rect 21324 13200 21330 13252
rect 21358 13200 21364 13252
rect 21416 13240 21422 13252
rect 21416 13212 22094 13240
rect 21416 13200 21422 13212
rect 15344 13144 16252 13172
rect 15344 13132 15350 13144
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 21542 13172 21548 13184
rect 16356 13144 21548 13172
rect 16356 13132 16362 13144
rect 21542 13132 21548 13144
rect 21600 13132 21606 13184
rect 22066 13172 22094 13212
rect 22186 13200 22192 13252
rect 22244 13200 22250 13252
rect 22646 13200 22652 13252
rect 22704 13200 22710 13252
rect 23566 13200 23572 13252
rect 23624 13240 23630 13252
rect 24949 13243 25007 13249
rect 24949 13240 24961 13243
rect 23624 13212 24961 13240
rect 23624 13200 23630 13212
rect 24949 13209 24961 13212
rect 24995 13209 25007 13243
rect 24949 13203 25007 13209
rect 23661 13175 23719 13181
rect 23661 13172 23673 13175
rect 22066 13144 23673 13172
rect 23661 13141 23673 13144
rect 23707 13141 23719 13175
rect 23661 13135 23719 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 14182 12968 14188 12980
rect 12912 12940 14188 12968
rect 12912 12841 12940 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14642 12928 14648 12980
rect 14700 12928 14706 12980
rect 19426 12968 19432 12980
rect 18524 12940 19432 12968
rect 13170 12860 13176 12912
rect 13228 12860 13234 12912
rect 13630 12860 13636 12912
rect 13688 12860 13694 12912
rect 16669 12903 16727 12909
rect 16669 12869 16681 12903
rect 16715 12900 16727 12903
rect 18322 12900 18328 12912
rect 16715 12872 18328 12900
rect 16715 12869 16727 12872
rect 16669 12863 16727 12869
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 17862 12832 17868 12844
rect 15151 12804 17868 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 18524 12841 18552 12940
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19794 12928 19800 12980
rect 19852 12968 19858 12980
rect 20809 12971 20867 12977
rect 20809 12968 20821 12971
rect 19852 12940 20821 12968
rect 19852 12928 19858 12940
rect 20809 12937 20821 12940
rect 20855 12937 20867 12971
rect 20809 12931 20867 12937
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 23753 12971 23811 12977
rect 23753 12968 23765 12971
rect 22244 12940 23765 12968
rect 22244 12928 22250 12940
rect 23753 12937 23765 12940
rect 23799 12968 23811 12971
rect 25130 12968 25136 12980
rect 23799 12940 25136 12968
rect 23799 12937 23811 12940
rect 23753 12931 23811 12937
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 18782 12860 18788 12912
rect 18840 12860 18846 12912
rect 20070 12900 20076 12912
rect 20010 12872 20076 12900
rect 20070 12860 20076 12872
rect 20128 12900 20134 12912
rect 21266 12900 21272 12912
rect 20128 12872 21272 12900
rect 20128 12860 20134 12872
rect 21266 12860 21272 12872
rect 21324 12860 21330 12912
rect 22922 12860 22928 12912
rect 22980 12860 22986 12912
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12801 18567 12835
rect 18509 12795 18567 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 15381 12767 15439 12773
rect 15381 12733 15393 12767
rect 15427 12764 15439 12767
rect 18230 12764 18236 12776
rect 15427 12736 18236 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 20732 12764 20760 12795
rect 25038 12792 25044 12844
rect 25096 12792 25102 12844
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 18616 12736 20760 12764
rect 20824 12736 20913 12764
rect 18616 12640 18644 12736
rect 20824 12708 20852 12736
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 22281 12767 22339 12773
rect 22281 12733 22293 12767
rect 22327 12764 22339 12767
rect 22327 12736 23428 12764
rect 22327 12733 22339 12736
rect 22281 12727 22339 12733
rect 20162 12656 20168 12708
rect 20220 12696 20226 12708
rect 20257 12699 20315 12705
rect 20257 12696 20269 12699
rect 20220 12668 20269 12696
rect 20220 12656 20226 12668
rect 20257 12665 20269 12668
rect 20303 12665 20315 12699
rect 20257 12659 20315 12665
rect 20806 12656 20812 12708
rect 20864 12656 20870 12708
rect 23400 12696 23428 12736
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 24397 12767 24455 12773
rect 24397 12764 24409 12767
rect 23532 12736 24409 12764
rect 23532 12724 23538 12736
rect 24397 12733 24409 12736
rect 24443 12733 24455 12767
rect 24397 12727 24455 12733
rect 23934 12696 23940 12708
rect 23400 12668 23940 12696
rect 23934 12656 23940 12668
rect 23992 12696 23998 12708
rect 24670 12696 24676 12708
rect 23992 12668 24676 12696
rect 23992 12656 23998 12668
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 17957 12631 18015 12637
rect 17957 12628 17969 12631
rect 17092 12600 17969 12628
rect 17092 12588 17098 12600
rect 17957 12597 17969 12600
rect 18003 12597 18015 12631
rect 17957 12591 18015 12597
rect 18598 12588 18604 12640
rect 18656 12588 18662 12640
rect 20346 12588 20352 12640
rect 20404 12588 20410 12640
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 23014 12628 23020 12640
rect 20496 12600 23020 12628
rect 20496 12588 20502 12600
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 18141 12427 18199 12433
rect 16724 12396 17172 12424
rect 16724 12384 16730 12396
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 15749 12291 15807 12297
rect 4212 12260 6914 12288
rect 4212 12248 4218 12260
rect 6886 12084 6914 12260
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 17034 12288 17040 12300
rect 15795 12260 17040 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 17144 12220 17172 12396
rect 18141 12393 18153 12427
rect 18187 12424 18199 12427
rect 18414 12424 18420 12436
rect 18187 12396 18420 12424
rect 18187 12393 18199 12396
rect 18141 12387 18199 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 19518 12384 19524 12436
rect 19576 12384 19582 12436
rect 19702 12433 19708 12436
rect 19692 12427 19708 12433
rect 19692 12393 19704 12427
rect 19760 12424 19766 12436
rect 21082 12424 21088 12436
rect 19760 12396 21088 12424
rect 19692 12387 19708 12393
rect 19702 12384 19708 12387
rect 19760 12384 19766 12396
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21358 12384 21364 12436
rect 21416 12424 21422 12436
rect 21726 12424 21732 12436
rect 21416 12396 21732 12424
rect 21416 12384 21422 12396
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 24029 12427 24087 12433
rect 24029 12393 24041 12427
rect 24075 12393 24087 12427
rect 24029 12387 24087 12393
rect 17218 12316 17224 12368
rect 17276 12356 17282 12368
rect 17497 12359 17555 12365
rect 17497 12356 17509 12359
rect 17276 12328 17509 12356
rect 17276 12316 17282 12328
rect 17497 12325 17509 12328
rect 17543 12356 17555 12359
rect 19536 12356 19564 12384
rect 17543 12328 19564 12356
rect 24044 12356 24072 12387
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24765 12427 24823 12433
rect 24765 12424 24777 12427
rect 24268 12396 24777 12424
rect 24268 12384 24274 12396
rect 24765 12393 24777 12396
rect 24811 12393 24823 12427
rect 24765 12387 24823 12393
rect 24670 12356 24676 12368
rect 24044 12328 24676 12356
rect 17543 12325 17555 12328
rect 17497 12319 17555 12325
rect 24670 12316 24676 12328
rect 24728 12316 24734 12368
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 20772 12260 21036 12288
rect 20772 12248 20778 12260
rect 18322 12220 18328 12232
rect 17144 12206 18328 12220
rect 17158 12192 18328 12206
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 19426 12180 19432 12232
rect 19484 12180 19490 12232
rect 16022 12112 16028 12164
rect 16080 12112 16086 12164
rect 18693 12155 18751 12161
rect 18693 12152 18705 12155
rect 17328 12124 18705 12152
rect 17328 12084 17356 12124
rect 18693 12121 18705 12124
rect 18739 12121 18751 12155
rect 18693 12115 18751 12121
rect 18877 12155 18935 12161
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 19334 12152 19340 12164
rect 18923 12124 19340 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 20162 12112 20168 12164
rect 20220 12112 20226 12164
rect 21008 12152 21036 12260
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21821 12291 21879 12297
rect 21821 12288 21833 12291
rect 21140 12260 21833 12288
rect 21140 12248 21146 12260
rect 21821 12257 21833 12260
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 24026 12288 24032 12300
rect 22603 12260 24032 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 22002 12220 22008 12232
rect 21232 12192 22008 12220
rect 21232 12180 21238 12192
rect 22002 12180 22008 12192
rect 22060 12220 22066 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22060 12192 22293 12220
rect 22060 12180 22066 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 21008 12124 21741 12152
rect 21729 12121 21741 12124
rect 21775 12121 21787 12155
rect 21729 12115 21787 12121
rect 22646 12112 22652 12164
rect 22704 12152 22710 12164
rect 22704 12124 23046 12152
rect 22704 12112 22710 12124
rect 6886 12056 17356 12084
rect 19610 12044 19616 12096
rect 19668 12084 19674 12096
rect 21082 12084 21088 12096
rect 19668 12056 21088 12084
rect 19668 12044 19674 12056
rect 21082 12044 21088 12056
rect 21140 12084 21146 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 21140 12056 21189 12084
rect 21140 12044 21146 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 21177 12047 21235 12053
rect 21269 12087 21327 12093
rect 21269 12053 21281 12087
rect 21315 12084 21327 12087
rect 21450 12084 21456 12096
rect 21315 12056 21456 12084
rect 21315 12053 21327 12056
rect 21269 12047 21327 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 21634 12044 21640 12096
rect 21692 12044 21698 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 14458 11840 14464 11892
rect 14516 11840 14522 11892
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 15838 11840 15844 11892
rect 15896 11840 15902 11892
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 15988 11852 16129 11880
rect 15988 11840 15994 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 16117 11843 16175 11849
rect 19153 11883 19211 11889
rect 19153 11849 19165 11883
rect 19199 11880 19211 11883
rect 19242 11880 19248 11892
rect 19199 11852 19248 11880
rect 19199 11849 19211 11852
rect 19153 11843 19211 11849
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 21174 11880 21180 11892
rect 19352 11852 21180 11880
rect 14001 11815 14059 11821
rect 14001 11781 14013 11815
rect 14047 11812 14059 11815
rect 16574 11812 16580 11824
rect 14047 11784 16580 11812
rect 14047 11781 14059 11784
rect 14001 11775 14059 11781
rect 14660 11753 14688 11784
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 17034 11812 17040 11824
rect 16868 11784 17040 11812
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15838 11744 15844 11756
rect 15335 11716 15844 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16298 11704 16304 11756
rect 16356 11704 16362 11756
rect 16868 11753 16896 11784
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 17129 11815 17187 11821
rect 17129 11781 17141 11815
rect 17175 11812 17187 11815
rect 17218 11812 17224 11824
rect 17175 11784 17224 11812
rect 17175 11781 17187 11784
rect 17129 11775 17187 11781
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 18138 11772 18144 11824
rect 18196 11772 18202 11824
rect 19352 11753 19380 11852
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 19610 11772 19616 11824
rect 19668 11772 19674 11824
rect 20070 11772 20076 11824
rect 20128 11772 20134 11824
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 21634 11704 21640 11756
rect 21692 11744 21698 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21692 11716 22017 11744
rect 21692 11704 21698 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 20070 11676 20076 11688
rect 14608 11648 20076 11676
rect 14608 11636 14614 11648
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 21085 11679 21143 11685
rect 21085 11676 21097 11679
rect 20312 11648 21097 11676
rect 20312 11636 20318 11648
rect 21085 11645 21097 11648
rect 21131 11676 21143 11679
rect 21542 11676 21548 11688
rect 21131 11648 21548 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 21910 11636 21916 11688
rect 21968 11676 21974 11688
rect 22112 11676 22140 11707
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23532 11716 23949 11744
rect 23532 11704 23538 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 21968 11648 22140 11676
rect 21968 11636 21974 11648
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 16850 11608 16856 11620
rect 14332 11580 16856 11608
rect 14332 11568 14338 11580
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 17678 11500 17684 11552
rect 17736 11540 17742 11552
rect 18601 11543 18659 11549
rect 18601 11540 18613 11543
rect 17736 11512 18613 11540
rect 17736 11500 17742 11512
rect 18601 11509 18613 11512
rect 18647 11540 18659 11543
rect 20622 11540 20628 11552
rect 18647 11512 20628 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 21082 11500 21088 11552
rect 21140 11540 21146 11552
rect 24578 11540 24584 11552
rect 21140 11512 24584 11540
rect 21140 11500 21146 11512
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 6604 11308 12434 11336
rect 6604 11296 6610 11308
rect 12406 11268 12434 11308
rect 16390 11296 16396 11348
rect 16448 11336 16454 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 16448 11308 16497 11336
rect 16448 11296 16454 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 16592 11308 20024 11336
rect 16592 11268 16620 11308
rect 12406 11240 16620 11268
rect 18877 11271 18935 11277
rect 18877 11237 18889 11271
rect 18923 11268 18935 11271
rect 19702 11268 19708 11280
rect 18923 11240 19708 11268
rect 18923 11237 18935 11240
rect 18877 11231 18935 11237
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 19426 11200 19432 11212
rect 17175 11172 19432 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 16025 11135 16083 11141
rect 16025 11101 16037 11135
rect 16071 11132 16083 11135
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16071 11104 16681 11132
rect 16071 11101 16083 11104
rect 16025 11095 16083 11101
rect 16669 11101 16681 11104
rect 16715 11132 16727 11135
rect 16942 11132 16948 11144
rect 16715 11104 16948 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 19996 11141 20024 11308
rect 20990 11296 20996 11348
rect 21048 11336 21054 11348
rect 21821 11339 21879 11345
rect 21821 11336 21833 11339
rect 21048 11308 21833 11336
rect 21048 11296 21054 11308
rect 21821 11305 21833 11308
rect 21867 11305 21879 11339
rect 21821 11299 21879 11305
rect 22002 11296 22008 11348
rect 22060 11336 22066 11348
rect 23934 11336 23940 11348
rect 22060 11308 23940 11336
rect 22060 11296 22066 11308
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 24578 11296 24584 11348
rect 24636 11296 24642 11348
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11268 21235 11271
rect 24026 11268 24032 11280
rect 21223 11240 24032 11268
rect 21223 11237 21235 11240
rect 21177 11231 21235 11237
rect 24026 11228 24032 11240
rect 24084 11228 24090 11280
rect 20070 11160 20076 11212
rect 20128 11160 20134 11212
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 23845 11203 23903 11209
rect 20220 11172 22692 11200
rect 20220 11160 20226 11172
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11101 20039 11135
rect 20088 11132 20116 11160
rect 20088 11104 21220 11132
rect 19981 11095 20039 11101
rect 17405 11067 17463 11073
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 17678 11064 17684 11076
rect 17451 11036 17684 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 17678 11024 17684 11036
rect 17736 11024 17742 11076
rect 18138 11024 18144 11076
rect 18196 11024 18202 11076
rect 20165 11067 20223 11073
rect 20165 11033 20177 11067
rect 20211 11064 20223 11067
rect 20622 11064 20628 11076
rect 20211 11036 20628 11064
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 21192 11064 21220 11104
rect 21266 11092 21272 11144
rect 21324 11132 21330 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 21324 11104 21373 11132
rect 21324 11092 21330 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21818 11092 21824 11144
rect 21876 11132 21882 11144
rect 22664 11141 22692 11172
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24946 11200 24952 11212
rect 23891 11172 24952 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 22005 11135 22063 11141
rect 22005 11132 22017 11135
rect 21876 11104 22017 11132
rect 21876 11092 21882 11104
rect 22005 11101 22017 11104
rect 22051 11101 22063 11135
rect 22005 11095 22063 11101
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 24394 11092 24400 11144
rect 24452 11132 24458 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 24452 11104 24777 11132
rect 24452 11092 24458 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 21192 11036 21680 11064
rect 18414 10956 18420 11008
rect 18472 10996 18478 11008
rect 18874 10996 18880 11008
rect 18472 10968 18880 10996
rect 18472 10956 18478 10968
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 21652 10996 21680 11036
rect 21726 11024 21732 11076
rect 21784 11064 21790 11076
rect 23290 11064 23296 11076
rect 21784 11036 23296 11064
rect 21784 11024 21790 11036
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 22002 10996 22008 11008
rect 21652 10968 22008 10996
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 17313 10795 17371 10801
rect 17313 10792 17325 10795
rect 16816 10764 17325 10792
rect 16816 10752 16822 10764
rect 17313 10761 17325 10764
rect 17359 10761 17371 10795
rect 17313 10755 17371 10761
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 18506 10792 18512 10804
rect 17727 10764 18512 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 18932 10764 22094 10792
rect 18932 10752 18938 10764
rect 17221 10727 17279 10733
rect 17221 10693 17233 10727
rect 17267 10724 17279 10727
rect 17586 10724 17592 10736
rect 17267 10696 17592 10724
rect 17267 10693 17279 10696
rect 17221 10687 17279 10693
rect 17586 10684 17592 10696
rect 17644 10724 17650 10736
rect 17644 10696 17908 10724
rect 17644 10684 17650 10696
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 15197 10659 15255 10665
rect 15197 10656 15209 10659
rect 10284 10628 15209 10656
rect 10284 10616 10290 10628
rect 15197 10625 15209 10628
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 17368 10628 17509 10656
rect 17368 10616 17374 10628
rect 17497 10625 17509 10628
rect 17543 10656 17555 10659
rect 17770 10656 17776 10668
rect 17543 10628 17776 10656
rect 17543 10625 17555 10628
rect 17497 10619 17555 10625
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 17880 10665 17908 10696
rect 17954 10684 17960 10736
rect 18012 10724 18018 10736
rect 20806 10724 20812 10736
rect 18012 10696 20812 10724
rect 18012 10684 18018 10696
rect 20806 10684 20812 10696
rect 20864 10684 20870 10736
rect 22066 10724 22094 10764
rect 23293 10727 23351 10733
rect 22066 10696 22140 10724
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 18598 10616 18604 10668
rect 18656 10616 18662 10668
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10656 19027 10659
rect 19242 10656 19248 10668
rect 19015 10628 19248 10656
rect 19015 10625 19027 10628
rect 18969 10619 19027 10625
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 19794 10656 19800 10668
rect 19659 10628 19800 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 19794 10616 19800 10628
rect 19852 10616 19858 10668
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10656 20315 10659
rect 20530 10656 20536 10668
rect 20303 10628 20536 10656
rect 20303 10625 20315 10628
rect 20257 10619 20315 10625
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 20898 10616 20904 10668
rect 20956 10616 20962 10668
rect 22112 10665 22140 10696
rect 23293 10693 23305 10727
rect 23339 10724 23351 10727
rect 24854 10724 24860 10736
rect 23339 10696 24860 10724
rect 23339 10693 23351 10696
rect 23293 10687 23351 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10588 15531 10591
rect 20162 10588 20168 10600
rect 15519 10560 20168 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 24670 10548 24676 10600
rect 24728 10548 24734 10600
rect 19978 10480 19984 10532
rect 20036 10520 20042 10532
rect 25130 10520 25136 10532
rect 20036 10492 25136 10520
rect 20036 10480 20042 10492
rect 25130 10480 25136 10492
rect 25188 10480 25194 10532
rect 19426 10412 19432 10464
rect 19484 10412 19490 10464
rect 20073 10455 20131 10461
rect 20073 10421 20085 10455
rect 20119 10452 20131 10455
rect 20162 10452 20168 10464
rect 20119 10424 20168 10452
rect 20119 10421 20131 10424
rect 20073 10415 20131 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 20717 10455 20775 10461
rect 20717 10421 20729 10455
rect 20763 10452 20775 10455
rect 21358 10452 21364 10464
rect 20763 10424 21364 10452
rect 20763 10421 20775 10424
rect 20717 10415 20775 10421
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22738 10452 22744 10464
rect 22336 10424 22744 10452
rect 22336 10412 22342 10424
rect 22738 10412 22744 10424
rect 22796 10412 22802 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 17310 10208 17316 10260
rect 17368 10208 17374 10260
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 17494 10248 17500 10260
rect 17451 10220 17500 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 19429 10251 19487 10257
rect 19429 10217 19441 10251
rect 19475 10248 19487 10251
rect 19518 10248 19524 10260
rect 19475 10220 19524 10248
rect 19475 10217 19487 10220
rect 19429 10211 19487 10217
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 23845 10251 23903 10257
rect 23845 10248 23857 10251
rect 21100 10220 23857 10248
rect 20714 10180 20720 10192
rect 17604 10152 20720 10180
rect 17604 10053 17632 10152
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 20254 10112 20260 10124
rect 18095 10084 20260 10112
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 21100 10112 21128 10220
rect 23845 10217 23857 10220
rect 23891 10217 23903 10251
rect 23845 10211 23903 10217
rect 24581 10183 24639 10189
rect 24581 10149 24593 10183
rect 24627 10149 24639 10183
rect 24581 10143 24639 10149
rect 20456 10084 21128 10112
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10044 19671 10047
rect 20070 10044 20076 10056
rect 19659 10016 20076 10044
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 18340 9976 18368 10007
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20456 10053 20484 10084
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 21232 10084 21281 10112
rect 21232 10072 21238 10084
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21542 10072 21548 10124
rect 21600 10072 21606 10124
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 24596 10112 24624 10143
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 22244 10084 24624 10112
rect 24688 10084 25145 10112
rect 22244 10072 22250 10084
rect 20441 10047 20499 10053
rect 20441 10013 20453 10047
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 20530 10004 20536 10056
rect 20588 10044 20594 10056
rect 20588 10016 20852 10044
rect 20588 10004 20594 10016
rect 20714 9976 20720 9988
rect 18340 9948 20720 9976
rect 20714 9936 20720 9948
rect 20772 9936 20778 9988
rect 20824 9976 20852 10016
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10044 24087 10047
rect 24118 10044 24124 10056
rect 24075 10016 24124 10044
rect 24075 10013 24087 10016
rect 24029 10007 24087 10013
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 21818 9976 21824 9988
rect 20824 9948 21824 9976
rect 21818 9936 21824 9948
rect 21876 9936 21882 9988
rect 23934 9976 23940 9988
rect 22940 9948 23940 9976
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9908 20315 9911
rect 22940 9908 22968 9948
rect 23934 9936 23940 9948
rect 23992 9936 23998 9988
rect 20303 9880 22968 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 23014 9868 23020 9920
rect 23072 9908 23078 9920
rect 24688 9908 24716 10084
rect 25133 10081 25145 10084
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25038 10044 25044 10056
rect 24995 10016 25044 10044
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 23072 9880 24716 9908
rect 25041 9911 25099 9917
rect 23072 9868 23078 9880
rect 25041 9877 25053 9911
rect 25087 9908 25099 9911
rect 25130 9908 25136 9920
rect 25087 9880 25136 9908
rect 25087 9877 25099 9880
rect 25041 9871 25099 9877
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 20070 9664 20076 9716
rect 20128 9704 20134 9716
rect 20530 9704 20536 9716
rect 20128 9676 20536 9704
rect 20128 9664 20134 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 20625 9707 20683 9713
rect 20625 9673 20637 9707
rect 20671 9673 20683 9707
rect 20625 9667 20683 9673
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 20640 9636 20668 9667
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 20772 9676 21680 9704
rect 20772 9664 20778 9676
rect 21652 9636 21680 9676
rect 21818 9664 21824 9716
rect 21876 9704 21882 9716
rect 23014 9704 23020 9716
rect 21876 9676 23020 9704
rect 21876 9664 21882 9676
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 17460 9608 20300 9636
rect 20640 9608 21404 9636
rect 21652 9608 22140 9636
rect 17460 9596 17466 9608
rect 17589 9571 17647 9577
rect 17589 9537 17601 9571
rect 17635 9568 17647 9571
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17635 9540 18245 9568
rect 17635 9537 17647 9540
rect 17589 9531 17647 9537
rect 18233 9537 18245 9540
rect 18279 9568 18291 9571
rect 18690 9568 18696 9580
rect 18279 9540 18696 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 18966 9568 18972 9580
rect 18923 9540 18972 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 20162 9528 20168 9580
rect 20220 9528 20226 9580
rect 20272 9568 20300 9608
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20272 9540 20821 9568
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 21376 9500 21404 9608
rect 22112 9577 22140 9608
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 22097 9571 22155 9577
rect 21499 9540 21772 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21744 9500 21772 9540
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 22370 9500 22376 9512
rect 21376 9472 21496 9500
rect 21744 9472 22376 9500
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 19337 9435 19395 9441
rect 19337 9432 19349 9435
rect 16172 9404 19349 9432
rect 16172 9392 16178 9404
rect 19337 9401 19349 9404
rect 19383 9401 19395 9435
rect 19337 9395 19395 9401
rect 19981 9435 20039 9441
rect 19981 9401 19993 9435
rect 20027 9432 20039 9435
rect 21468 9432 21496 9472
rect 22370 9460 22376 9472
rect 22428 9460 22434 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 24302 9432 24308 9444
rect 20027 9404 21404 9432
rect 21468 9404 24308 9432
rect 20027 9401 20039 9404
rect 19981 9395 20039 9401
rect 18046 9324 18052 9376
rect 18104 9324 18110 9376
rect 18690 9324 18696 9376
rect 18748 9324 18754 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20312 9336 21281 9364
rect 20312 9324 20318 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21376 9364 21404 9404
rect 24302 9392 24308 9404
rect 24360 9392 24366 9444
rect 23382 9364 23388 9376
rect 21376 9336 23388 9364
rect 21269 9327 21327 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 14366 9160 14372 9172
rect 11931 9132 14372 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 26050 9160 26056 9172
rect 19576 9132 26056 9160
rect 19576 9120 19582 9132
rect 26050 9120 26056 9132
rect 26108 9120 26114 9172
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 21361 9095 21419 9101
rect 21361 9092 21373 9095
rect 16908 9064 21373 9092
rect 16908 9052 16914 9064
rect 21361 9061 21373 9064
rect 21407 9061 21419 9095
rect 25682 9092 25688 9104
rect 21361 9055 21419 9061
rect 22066 9064 25688 9092
rect 10134 8984 10140 9036
rect 10192 8984 10198 9036
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 18748 8996 19441 9024
rect 18748 8984 18754 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20806 8956 20812 8968
rect 19751 8928 20812 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20806 8916 20812 8928
rect 20864 8916 20870 8968
rect 20901 8959 20959 8965
rect 20901 8925 20913 8959
rect 20947 8925 20959 8959
rect 20901 8919 20959 8925
rect 21545 8959 21603 8965
rect 21545 8925 21557 8959
rect 21591 8956 21603 8959
rect 22066 8956 22094 9064
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24946 9024 24952 9036
rect 23891 8996 24952 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24946 8984 24952 8996
rect 25004 8984 25010 9036
rect 21591 8928 22094 8956
rect 22189 8959 22247 8965
rect 21591 8925 21603 8928
rect 21545 8919 21603 8925
rect 22189 8925 22201 8959
rect 22235 8956 22247 8959
rect 22554 8956 22560 8968
rect 22235 8928 22560 8956
rect 22235 8925 22247 8928
rect 22189 8919 22247 8925
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 10413 8891 10471 8897
rect 10413 8888 10425 8891
rect 6880 8860 10425 8888
rect 6880 8848 6886 8860
rect 10413 8857 10425 8860
rect 10459 8857 10471 8891
rect 12342 8888 12348 8900
rect 11638 8860 12348 8888
rect 10413 8851 10471 8857
rect 12342 8848 12348 8860
rect 12400 8848 12406 8900
rect 20916 8888 20944 8919
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 24394 8888 24400 8900
rect 20916 8860 24400 8888
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 24673 8891 24731 8897
rect 24673 8857 24685 8891
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 24857 8891 24915 8897
rect 24857 8857 24869 8891
rect 24903 8888 24915 8891
rect 25130 8888 25136 8900
rect 24903 8860 25136 8888
rect 24903 8857 24915 8860
rect 24857 8851 24915 8857
rect 20714 8780 20720 8832
rect 20772 8780 20778 8832
rect 22005 8823 22063 8829
rect 22005 8789 22017 8823
rect 22051 8820 22063 8823
rect 24688 8820 24716 8851
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 22051 8792 24716 8820
rect 22051 8789 22063 8792
rect 22005 8783 22063 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 14792 8588 19993 8616
rect 14792 8576 14798 8588
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 19981 8579 20039 8585
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 23474 8616 23480 8628
rect 21315 8588 23480 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 20346 8508 20352 8560
rect 20404 8548 20410 8560
rect 20404 8520 20576 8548
rect 20404 8508 20410 8520
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8480 20223 8483
rect 20438 8480 20444 8492
rect 20211 8452 20444 8480
rect 20211 8449 20223 8452
rect 20165 8443 20223 8449
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20548 8480 20576 8520
rect 20714 8508 20720 8560
rect 20772 8548 20778 8560
rect 23293 8551 23351 8557
rect 20772 8520 22416 8548
rect 20772 8508 20778 8520
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20548 8452 20821 8480
rect 20809 8449 20821 8452
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8480 21511 8483
rect 21726 8480 21732 8492
rect 21499 8452 21732 8480
rect 21499 8449 21511 8452
rect 21453 8443 21511 8449
rect 21726 8440 21732 8452
rect 21784 8440 21790 8492
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22388 8480 22416 8520
rect 23293 8517 23305 8551
rect 23339 8548 23351 8551
rect 24854 8548 24860 8560
rect 23339 8520 24860 8548
rect 23339 8517 23351 8520
rect 23293 8511 23351 8517
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 22388 8452 23949 8480
rect 22281 8443 22339 8449
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 25222 8480 25228 8492
rect 23937 8443 23995 8449
rect 24044 8452 25228 8480
rect 22296 8412 22324 8443
rect 24044 8412 24072 8452
rect 25222 8440 25228 8452
rect 25280 8440 25286 8492
rect 22296 8384 24072 8412
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 20625 8347 20683 8353
rect 20625 8313 20637 8347
rect 20671 8344 20683 8347
rect 24026 8344 24032 8356
rect 20671 8316 24032 8344
rect 20671 8313 20683 8316
rect 20625 8307 20683 8313
rect 24026 8304 24032 8316
rect 24084 8304 24090 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 20717 8075 20775 8081
rect 20717 8041 20729 8075
rect 20763 8072 20775 8075
rect 22646 8072 22652 8084
rect 20763 8044 22652 8072
rect 20763 8041 20775 8044
rect 20717 8035 20775 8041
rect 22646 8032 22652 8044
rect 22704 8032 22710 8084
rect 24394 8032 24400 8084
rect 24452 8072 24458 8084
rect 24581 8075 24639 8081
rect 24581 8072 24593 8075
rect 24452 8044 24593 8072
rect 24452 8032 24458 8044
rect 24581 8041 24593 8044
rect 24627 8041 24639 8075
rect 24581 8035 24639 8041
rect 21361 8007 21419 8013
rect 21361 7973 21373 8007
rect 21407 8004 21419 8007
rect 21910 8004 21916 8016
rect 21407 7976 21916 8004
rect 21407 7973 21419 7976
rect 21361 7967 21419 7973
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 22189 8007 22247 8013
rect 22189 7973 22201 8007
rect 22235 8004 22247 8007
rect 23566 8004 23572 8016
rect 22235 7976 23572 8004
rect 22235 7973 22247 7976
rect 22189 7967 22247 7973
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 23845 7939 23903 7945
rect 21692 7908 23428 7936
rect 21692 7896 21698 7908
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 19484 7840 20913 7868
rect 19484 7828 19490 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21542 7828 21548 7880
rect 21600 7828 21606 7880
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 23400 7868 23428 7908
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24946 7936 24952 7948
rect 23891 7908 24952 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24946 7896 24952 7908
rect 25004 7896 25010 7948
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 23400 7840 24777 7868
rect 22833 7831 22891 7837
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 22848 7800 22876 7831
rect 24854 7800 24860 7812
rect 22848 7772 24860 7800
rect 24854 7760 24860 7772
rect 24912 7760 24918 7812
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 25406 7528 25412 7540
rect 23216 7500 25412 7528
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 23216 7392 23244 7500
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 23293 7463 23351 7469
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 22327 7364 23244 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 23382 7352 23388 7404
rect 23440 7392 23446 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23440 7364 23949 7392
rect 23440 7352 23446 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24670 7284 24676 7336
rect 24728 7284 24734 7336
rect 20809 7259 20867 7265
rect 20809 7225 20821 7259
rect 20855 7256 20867 7259
rect 25038 7256 25044 7268
rect 20855 7228 25044 7256
rect 20855 7225 20867 7228
rect 20809 7219 20867 7225
rect 25038 7216 25044 7228
rect 25096 7216 25102 7268
rect 21269 7191 21327 7197
rect 21269 7157 21281 7191
rect 21315 7188 21327 7191
rect 22738 7188 22744 7200
rect 21315 7160 22744 7188
rect 21315 7157 21327 7160
rect 21269 7151 21327 7157
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 21361 6919 21419 6925
rect 21361 6885 21373 6919
rect 21407 6885 21419 6919
rect 21361 6879 21419 6885
rect 21376 6848 21404 6879
rect 23845 6851 23903 6857
rect 21376 6820 22692 6848
rect 21358 6740 21364 6792
rect 21416 6780 21422 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 21416 6752 21557 6780
rect 21416 6740 21422 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6780 22247 6783
rect 22278 6780 22284 6792
rect 22235 6752 22284 6780
rect 22235 6749 22247 6752
rect 22189 6743 22247 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 22664 6789 22692 6820
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24854 6848 24860 6860
rect 23891 6820 24860 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 24302 6740 24308 6792
rect 24360 6780 24366 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 24360 6752 24685 6780
rect 24360 6740 24366 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 11606 6672 11612 6724
rect 11664 6712 11670 6724
rect 24857 6715 24915 6721
rect 11664 6684 22048 6712
rect 11664 6672 11670 6684
rect 22020 6653 22048 6684
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25038 6712 25044 6724
rect 24903 6684 25044 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 22005 6647 22063 6653
rect 22005 6613 22017 6647
rect 22051 6613 22063 6647
rect 22005 6607 22063 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 25130 6440 25136 6452
rect 22296 6412 25136 6440
rect 22296 6313 22324 6412
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 24854 6372 24860 6384
rect 23339 6344 24860 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6304 24179 6307
rect 24486 6304 24492 6316
rect 24167 6276 24492 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 24486 6264 24492 6276
rect 24544 6264 24550 6316
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 22005 5831 22063 5837
rect 22005 5797 22017 5831
rect 22051 5828 22063 5831
rect 23290 5828 23296 5840
rect 22051 5800 23296 5828
rect 22051 5797 22063 5800
rect 22005 5791 22063 5797
rect 23290 5788 23296 5800
rect 23348 5788 23354 5840
rect 22186 5652 22192 5704
rect 22244 5652 22250 5704
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 22848 5556 22876 5655
rect 24118 5652 24124 5704
rect 24176 5692 24182 5704
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 24176 5664 24869 5692
rect 24176 5652 24182 5664
rect 24857 5661 24869 5664
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 24946 5624 24952 5636
rect 23891 5596 24952 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 22848 5528 24685 5556
rect 24673 5525 24685 5528
rect 24719 5525 24731 5559
rect 24673 5519 24731 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 20806 5244 20812 5296
rect 20864 5284 20870 5296
rect 23293 5287 23351 5293
rect 20864 5256 22232 5284
rect 20864 5244 20870 5256
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 22204 5216 22232 5256
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24854 5284 24860 5296
rect 23339 5256 24860 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 22204 5188 23949 5216
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 22462 4564 22468 4616
rect 22520 4604 22526 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22520 4576 22661 4604
rect 22520 4564 22526 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 24026 4564 24032 4616
rect 24084 4604 24090 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 24084 4576 24869 4604
rect 24084 4564 24090 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24946 4536 24952 4548
rect 23891 4508 24952 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 24670 4428 24676 4480
rect 24728 4428 24734 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 21174 4128 21180 4140
rect 20303 4100 21180 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 21174 4088 21180 4100
rect 21232 4088 21238 4140
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 22327 4100 22784 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 20162 4060 20168 4072
rect 17184 4032 20168 4060
rect 17184 4020 17190 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 22186 4060 22192 4072
rect 21315 4032 22192 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22186 4020 22192 4032
rect 22244 4020 22250 4072
rect 22756 3924 22784 4100
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 22888 4100 23949 4128
rect 22888 4088 22894 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 23308 3964 24952 3992
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 25038 3924 25044 3936
rect 22756 3896 25044 3924
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 22796 3556 24900 3584
rect 22796 3544 22802 3556
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20680 3488 20821 3516
rect 20680 3476 20686 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 24670 3516 24676 3528
rect 22879 3488 24676 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24872 3525 24900 3556
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24946 3448 24952 3460
rect 23891 3420 24952 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 22278 3340 22284 3392
rect 22336 3380 22342 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 22336 3352 24685 3380
rect 22336 3340 22342 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 24673 3343 24731 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 23293 3111 23351 3117
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 25130 3068 25136 3120
rect 25188 3068 25194 3120
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 18782 3040 18788 3052
rect 18463 3012 18788 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 19392 3012 20085 3040
rect 19392 3000 19398 3012
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 22278 3000 22284 3052
rect 22336 3000 22342 3052
rect 23842 3000 23848 3052
rect 23900 3040 23906 3052
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23900 3012 23949 3040
rect 23900 3000 23906 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19518 2972 19524 2984
rect 19475 2944 19524 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 25038 2972 25044 2984
rect 21315 2944 25044 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6822 2592 6828 2644
rect 6880 2592 6886 2644
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 23382 2496 23388 2508
rect 21315 2468 23388 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6788 2400 7021 2428
rect 6788 2388 6794 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 19518 2320 19524 2372
rect 19576 2360 19582 2372
rect 22094 2360 22100 2372
rect 19576 2332 22100 2360
rect 19576 2320 19582 2332
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 22848 2292 22876 2391
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 23348 2400 24777 2428
rect 23348 2388 23354 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 22848 2264 24593 2292
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 3056 26392 3108 26444
rect 3332 26392 3384 26444
rect 2228 26324 2280 26376
rect 22192 26324 22244 26376
rect 21456 26256 21508 26308
rect 5264 26188 5316 26240
rect 10232 24896 10284 24948
rect 20720 24896 20772 24948
rect 18512 24828 18564 24880
rect 18788 24828 18840 24880
rect 11520 24760 11572 24812
rect 13452 24760 13504 24812
rect 14188 24760 14240 24812
rect 23388 24760 23440 24812
rect 6552 24692 6604 24744
rect 13912 24692 13964 24744
rect 16580 24692 16632 24744
rect 21088 24692 21140 24744
rect 4896 24624 4948 24676
rect 14740 24624 14792 24676
rect 16028 24624 16080 24676
rect 22008 24624 22060 24676
rect 4804 24556 4856 24608
rect 15476 24556 15528 24608
rect 16396 24556 16448 24608
rect 24216 24556 24268 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 12716 24284 12768 24336
rect 18512 24352 18564 24404
rect 6460 24216 6512 24268
rect 3884 24148 3936 24200
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 5448 24148 5500 24200
rect 7012 24148 7064 24200
rect 9680 24216 9732 24268
rect 10968 24259 11020 24268
rect 10968 24225 10977 24259
rect 10977 24225 11011 24259
rect 11011 24225 11020 24259
rect 10968 24216 11020 24225
rect 12440 24216 12492 24268
rect 13912 24216 13964 24268
rect 16120 24216 16172 24268
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 19800 24284 19852 24336
rect 8668 24080 8720 24132
rect 9588 24148 9640 24200
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 13728 24148 13780 24200
rect 14280 24080 14332 24132
rect 14372 24123 14424 24132
rect 14372 24089 14381 24123
rect 14381 24089 14415 24123
rect 14415 24089 14424 24123
rect 14372 24080 14424 24089
rect 14556 24080 14608 24132
rect 3700 24012 3752 24064
rect 7104 24012 7156 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 9680 24012 9732 24064
rect 16580 24012 16632 24064
rect 16764 24123 16816 24132
rect 16764 24089 16773 24123
rect 16773 24089 16807 24123
rect 16807 24089 16816 24123
rect 16764 24080 16816 24089
rect 19156 24216 19208 24268
rect 21824 24352 21876 24404
rect 20720 24284 20772 24336
rect 21916 24216 21968 24268
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 20444 24148 20496 24200
rect 21088 24191 21140 24200
rect 21088 24157 21097 24191
rect 21097 24157 21131 24191
rect 21131 24157 21140 24191
rect 21088 24148 21140 24157
rect 21364 24148 21416 24200
rect 24492 24148 24544 24200
rect 17500 24080 17552 24132
rect 22560 24080 22612 24132
rect 22836 24123 22888 24132
rect 22836 24089 22845 24123
rect 22845 24089 22879 24123
rect 22879 24089 22888 24123
rect 22836 24080 22888 24089
rect 23848 24080 23900 24132
rect 19340 24012 19392 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 19892 24055 19944 24064
rect 19892 24021 19901 24055
rect 19901 24021 19935 24055
rect 19935 24021 19944 24055
rect 19892 24012 19944 24021
rect 23940 24012 23992 24064
rect 25044 24055 25096 24064
rect 25044 24021 25053 24055
rect 25053 24021 25087 24055
rect 25087 24021 25096 24055
rect 25044 24012 25096 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 4160 23808 4212 23860
rect 5080 23740 5132 23792
rect 7564 23740 7616 23792
rect 10140 23740 10192 23792
rect 10876 23783 10928 23792
rect 10876 23749 10885 23783
rect 10885 23749 10919 23783
rect 10919 23749 10928 23783
rect 10876 23740 10928 23749
rect 11888 23808 11940 23860
rect 14280 23808 14332 23860
rect 25044 23808 25096 23860
rect 940 23672 992 23724
rect 4896 23672 4948 23724
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 6736 23604 6788 23656
rect 7288 23672 7340 23724
rect 8392 23672 8444 23724
rect 8484 23604 8536 23656
rect 4344 23536 4396 23588
rect 17132 23740 17184 23792
rect 18420 23740 18472 23792
rect 18696 23740 18748 23792
rect 14280 23672 14332 23724
rect 22468 23740 22520 23792
rect 22836 23740 22888 23792
rect 24768 23740 24820 23792
rect 12256 23604 12308 23656
rect 14556 23647 14608 23656
rect 14556 23613 14565 23647
rect 14565 23613 14599 23647
rect 14599 23613 14608 23647
rect 14556 23604 14608 23613
rect 6552 23468 6604 23520
rect 7012 23468 7064 23520
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 16028 23647 16080 23656
rect 16028 23613 16037 23647
rect 16037 23613 16071 23647
rect 16071 23613 16080 23647
rect 16028 23604 16080 23613
rect 16120 23604 16172 23656
rect 16304 23604 16356 23656
rect 17316 23647 17368 23656
rect 17316 23613 17325 23647
rect 17325 23613 17359 23647
rect 17359 23613 17368 23647
rect 17316 23604 17368 23613
rect 17500 23647 17552 23656
rect 17500 23613 17509 23647
rect 17509 23613 17543 23647
rect 17543 23613 17552 23647
rect 17500 23604 17552 23613
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 19156 23604 19208 23656
rect 21272 23604 21324 23656
rect 22100 23647 22152 23656
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 22468 23604 22520 23656
rect 23848 23647 23900 23656
rect 23848 23613 23857 23647
rect 23857 23613 23891 23647
rect 23891 23613 23900 23647
rect 23848 23604 23900 23613
rect 19248 23536 19300 23588
rect 19708 23536 19760 23588
rect 20168 23536 20220 23588
rect 18880 23468 18932 23520
rect 19616 23511 19668 23520
rect 19616 23477 19625 23511
rect 19625 23477 19659 23511
rect 19659 23477 19668 23511
rect 19616 23468 19668 23477
rect 19800 23468 19852 23520
rect 20352 23468 20404 23520
rect 25596 23536 25648 23588
rect 25228 23511 25280 23520
rect 25228 23477 25237 23511
rect 25237 23477 25271 23511
rect 25271 23477 25280 23511
rect 25228 23468 25280 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 4160 23264 4212 23316
rect 9680 23264 9732 23316
rect 9956 23264 10008 23316
rect 14924 23264 14976 23316
rect 16304 23264 16356 23316
rect 19156 23264 19208 23316
rect 5080 23196 5132 23248
rect 5356 23196 5408 23248
rect 4620 23128 4672 23180
rect 7656 23196 7708 23248
rect 3608 23060 3660 23112
rect 4344 23060 4396 23112
rect 5632 23060 5684 23112
rect 7380 23128 7432 23180
rect 9404 23196 9456 23248
rect 10140 23196 10192 23248
rect 13912 23196 13964 23248
rect 18512 23196 18564 23248
rect 8576 23128 8628 23180
rect 9772 23060 9824 23112
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 11612 23128 11664 23180
rect 13544 23128 13596 23180
rect 15936 23128 15988 23180
rect 17868 23128 17920 23180
rect 21456 23196 21508 23248
rect 22008 23264 22060 23316
rect 22284 23264 22336 23316
rect 24032 23264 24084 23316
rect 23204 23196 23256 23248
rect 24952 23196 25004 23248
rect 21824 23171 21876 23180
rect 21824 23137 21833 23171
rect 21833 23137 21867 23171
rect 21867 23137 21876 23171
rect 21824 23128 21876 23137
rect 22284 23128 22336 23180
rect 11704 23103 11756 23112
rect 11704 23069 11713 23103
rect 11713 23069 11747 23103
rect 11747 23069 11756 23103
rect 11704 23060 11756 23069
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 1952 22924 2004 22976
rect 4160 22924 4212 22976
rect 11704 22924 11756 22976
rect 15476 22992 15528 23044
rect 15660 22992 15712 23044
rect 14096 22924 14148 22976
rect 17224 22924 17276 22976
rect 17960 22992 18012 23044
rect 19248 22992 19300 23044
rect 19708 23035 19760 23044
rect 19708 23001 19717 23035
rect 19717 23001 19751 23035
rect 19751 23001 19760 23035
rect 19708 22992 19760 23001
rect 19984 22992 20036 23044
rect 17500 22924 17552 22976
rect 19524 22924 19576 22976
rect 19616 22924 19668 22976
rect 21916 22992 21968 23044
rect 21640 22924 21692 22976
rect 21732 22924 21784 22976
rect 22008 22924 22060 22976
rect 23112 22992 23164 23044
rect 24032 22992 24084 23044
rect 22836 22924 22888 22976
rect 23388 22924 23440 22976
rect 24860 22924 24912 22976
rect 25412 22924 25464 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 8576 22720 8628 22772
rect 9496 22720 9548 22772
rect 4252 22652 4304 22704
rect 4436 22652 4488 22704
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 940 22584 992 22636
rect 4528 22584 4580 22636
rect 5172 22584 5224 22636
rect 6644 22627 6696 22636
rect 6644 22593 6653 22627
rect 6653 22593 6687 22627
rect 6687 22593 6696 22627
rect 6644 22584 6696 22593
rect 6828 22584 6880 22636
rect 7748 22584 7800 22636
rect 9956 22652 10008 22704
rect 11336 22652 11388 22704
rect 12256 22652 12308 22704
rect 12624 22652 12676 22704
rect 11428 22584 11480 22636
rect 13360 22584 13412 22636
rect 9128 22516 9180 22568
rect 12164 22516 12216 22568
rect 12348 22516 12400 22568
rect 14556 22720 14608 22772
rect 15936 22763 15988 22772
rect 15936 22729 15945 22763
rect 15945 22729 15979 22763
rect 15979 22729 15988 22763
rect 15936 22720 15988 22729
rect 17040 22763 17092 22772
rect 17040 22729 17049 22763
rect 17049 22729 17083 22763
rect 17083 22729 17092 22763
rect 17040 22720 17092 22729
rect 17132 22720 17184 22772
rect 17408 22720 17460 22772
rect 18512 22720 18564 22772
rect 18880 22720 18932 22772
rect 19984 22720 20036 22772
rect 22008 22720 22060 22772
rect 22284 22720 22336 22772
rect 14096 22652 14148 22704
rect 14280 22652 14332 22704
rect 16488 22652 16540 22704
rect 19156 22652 19208 22704
rect 20260 22652 20312 22704
rect 20444 22652 20496 22704
rect 25228 22720 25280 22772
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 15108 22584 15160 22636
rect 15752 22584 15804 22636
rect 7012 22448 7064 22500
rect 11152 22491 11204 22500
rect 11152 22457 11161 22491
rect 11161 22457 11195 22491
rect 11195 22457 11204 22491
rect 11152 22448 11204 22457
rect 11888 22448 11940 22500
rect 6736 22423 6788 22432
rect 6736 22389 6745 22423
rect 6745 22389 6779 22423
rect 6779 22389 6788 22423
rect 6736 22380 6788 22389
rect 9312 22380 9364 22432
rect 12256 22380 12308 22432
rect 12624 22380 12676 22432
rect 15568 22516 15620 22568
rect 16856 22584 16908 22636
rect 16304 22516 16356 22568
rect 17224 22584 17276 22636
rect 18420 22584 18472 22636
rect 20536 22627 20588 22636
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 21824 22584 21876 22636
rect 24492 22627 24544 22636
rect 24492 22593 24501 22627
rect 24501 22593 24535 22627
rect 24535 22593 24544 22627
rect 24492 22584 24544 22593
rect 15844 22448 15896 22500
rect 16580 22448 16632 22500
rect 16856 22448 16908 22500
rect 17592 22448 17644 22500
rect 19432 22559 19484 22568
rect 19432 22525 19441 22559
rect 19441 22525 19475 22559
rect 19475 22525 19484 22559
rect 19432 22516 19484 22525
rect 19524 22516 19576 22568
rect 17868 22448 17920 22500
rect 18328 22448 18380 22500
rect 19800 22448 19852 22500
rect 19984 22448 20036 22500
rect 16396 22380 16448 22432
rect 16948 22380 17000 22432
rect 19524 22380 19576 22432
rect 20076 22380 20128 22432
rect 22284 22448 22336 22500
rect 22468 22559 22520 22568
rect 22468 22525 22477 22559
rect 22477 22525 22511 22559
rect 22511 22525 22520 22559
rect 22468 22516 22520 22525
rect 22836 22516 22888 22568
rect 22560 22448 22612 22500
rect 24676 22559 24728 22568
rect 24676 22525 24685 22559
rect 24685 22525 24719 22559
rect 24719 22525 24728 22559
rect 24676 22516 24728 22525
rect 20996 22380 21048 22432
rect 21732 22380 21784 22432
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 22192 22380 22244 22432
rect 23112 22380 23164 22432
rect 23664 22423 23716 22432
rect 23664 22389 23673 22423
rect 23673 22389 23707 22423
rect 23707 22389 23716 22423
rect 23664 22380 23716 22389
rect 25044 22380 25096 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 9772 22176 9824 22228
rect 13636 22176 13688 22228
rect 2044 22108 2096 22160
rect 2964 22108 3016 22160
rect 3608 22108 3660 22160
rect 10508 22108 10560 22160
rect 11888 22108 11940 22160
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8300 22083 8352 22092
rect 8300 22049 8309 22083
rect 8309 22049 8343 22083
rect 8343 22049 8352 22083
rect 8300 22040 8352 22049
rect 9128 22040 9180 22092
rect 3424 21972 3476 22024
rect 4528 21972 4580 22024
rect 4804 21972 4856 22024
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 7472 21972 7524 22024
rect 4528 21836 4580 21888
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 9864 21904 9916 21956
rect 7840 21836 7892 21888
rect 8852 21836 8904 21888
rect 10140 22015 10192 22024
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 12164 22040 12216 22092
rect 13268 22108 13320 22160
rect 13728 22108 13780 22160
rect 14004 22108 14056 22160
rect 14372 22108 14424 22160
rect 14740 22108 14792 22160
rect 15200 22040 15252 22092
rect 15476 22040 15528 22092
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 12440 21972 12492 22024
rect 13728 21972 13780 22024
rect 15016 21972 15068 22024
rect 15108 21972 15160 22024
rect 11336 21904 11388 21956
rect 14096 21904 14148 21956
rect 14648 21947 14700 21956
rect 14648 21913 14657 21947
rect 14657 21913 14691 21947
rect 14691 21913 14700 21947
rect 14648 21904 14700 21913
rect 15384 21947 15436 21956
rect 15384 21913 15393 21947
rect 15393 21913 15427 21947
rect 15427 21913 15436 21947
rect 15384 21904 15436 21913
rect 13452 21836 13504 21888
rect 16396 21972 16448 22024
rect 18604 22176 18656 22228
rect 18880 22176 18932 22228
rect 20812 22176 20864 22228
rect 21732 22176 21784 22228
rect 21916 22176 21968 22228
rect 17408 22040 17460 22092
rect 18512 22040 18564 22092
rect 22284 22108 22336 22160
rect 20076 22083 20128 22092
rect 20076 22049 20085 22083
rect 20085 22049 20119 22083
rect 20119 22049 20128 22083
rect 20076 22040 20128 22049
rect 22100 22040 22152 22092
rect 22376 22040 22428 22092
rect 23296 22108 23348 22160
rect 23480 22108 23532 22160
rect 24492 22108 24544 22160
rect 25136 22108 25188 22160
rect 25412 22040 25464 22092
rect 16120 21836 16172 21888
rect 16764 21836 16816 21888
rect 17868 21904 17920 21956
rect 18604 21947 18656 21956
rect 18604 21913 18613 21947
rect 18613 21913 18647 21947
rect 18647 21913 18656 21947
rect 18604 21904 18656 21913
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 23296 21972 23348 22024
rect 20996 21904 21048 21956
rect 21732 21904 21784 21956
rect 19708 21836 19760 21888
rect 21364 21836 21416 21888
rect 23480 21836 23532 21888
rect 23572 21836 23624 21888
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 25320 21836 25372 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 2780 21632 2832 21684
rect 6736 21564 6788 21616
rect 10876 21564 10928 21616
rect 11336 21564 11388 21616
rect 12072 21675 12124 21684
rect 12072 21641 12081 21675
rect 12081 21641 12115 21675
rect 12115 21641 12124 21675
rect 12072 21632 12124 21641
rect 12440 21675 12492 21684
rect 12440 21641 12449 21675
rect 12449 21641 12483 21675
rect 12483 21641 12492 21675
rect 12440 21632 12492 21641
rect 13268 21564 13320 21616
rect 14556 21632 14608 21684
rect 16028 21632 16080 21684
rect 17040 21632 17092 21684
rect 17408 21632 17460 21684
rect 17684 21632 17736 21684
rect 13820 21564 13872 21616
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 8576 21496 8628 21548
rect 12164 21496 12216 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 4988 21428 5040 21480
rect 7196 21428 7248 21480
rect 9128 21471 9180 21480
rect 9128 21437 9137 21471
rect 9137 21437 9171 21471
rect 9171 21437 9180 21471
rect 9128 21428 9180 21437
rect 11152 21428 11204 21480
rect 12532 21471 12584 21480
rect 12532 21437 12541 21471
rect 12541 21437 12575 21471
rect 12575 21437 12584 21471
rect 12532 21428 12584 21437
rect 12716 21428 12768 21480
rect 15016 21496 15068 21548
rect 15292 21496 15344 21548
rect 17408 21539 17460 21548
rect 17408 21505 17417 21539
rect 17417 21505 17451 21539
rect 17451 21505 17460 21539
rect 17408 21496 17460 21505
rect 17776 21496 17828 21548
rect 18788 21564 18840 21616
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 20260 21632 20312 21684
rect 23572 21632 23624 21684
rect 24032 21675 24084 21684
rect 24032 21641 24041 21675
rect 24041 21641 24075 21675
rect 24075 21641 24084 21675
rect 24032 21632 24084 21641
rect 25044 21675 25096 21684
rect 25044 21641 25053 21675
rect 25053 21641 25087 21675
rect 25087 21641 25096 21675
rect 25044 21632 25096 21641
rect 22652 21564 22704 21616
rect 23848 21564 23900 21616
rect 19616 21496 19668 21548
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 21364 21496 21416 21548
rect 25044 21496 25096 21548
rect 10416 21360 10468 21412
rect 15476 21428 15528 21480
rect 16028 21428 16080 21480
rect 17500 21428 17552 21480
rect 17684 21471 17736 21480
rect 17684 21437 17693 21471
rect 17693 21437 17727 21471
rect 17727 21437 17736 21471
rect 17684 21428 17736 21437
rect 18512 21471 18564 21480
rect 18512 21437 18521 21471
rect 18521 21437 18555 21471
rect 18555 21437 18564 21471
rect 18512 21428 18564 21437
rect 18880 21428 18932 21480
rect 21272 21428 21324 21480
rect 22100 21428 22152 21480
rect 10140 21292 10192 21344
rect 10692 21292 10744 21344
rect 10968 21292 11020 21344
rect 12440 21292 12492 21344
rect 12532 21292 12584 21344
rect 13728 21292 13780 21344
rect 14096 21292 14148 21344
rect 15016 21335 15068 21344
rect 15016 21301 15025 21335
rect 15025 21301 15059 21335
rect 15059 21301 15068 21335
rect 15016 21292 15068 21301
rect 15384 21360 15436 21412
rect 18052 21360 18104 21412
rect 22560 21428 22612 21480
rect 22652 21428 22704 21480
rect 16672 21292 16724 21344
rect 23756 21360 23808 21412
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 20996 21292 21048 21344
rect 22008 21292 22060 21344
rect 22376 21292 22428 21344
rect 23664 21292 23716 21344
rect 25688 21292 25740 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2044 21088 2096 21140
rect 7748 21088 7800 21140
rect 2780 21020 2832 21072
rect 6920 21020 6972 21072
rect 7012 21020 7064 21072
rect 4160 20952 4212 21004
rect 5724 20884 5776 20936
rect 6552 20884 6604 20936
rect 7656 20884 7708 20936
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 12440 21020 12492 21072
rect 13636 21088 13688 21140
rect 16856 21131 16908 21140
rect 16856 21097 16865 21131
rect 16865 21097 16899 21131
rect 16899 21097 16908 21131
rect 16856 21088 16908 21097
rect 16948 21088 17000 21140
rect 10692 20952 10744 21004
rect 14280 21063 14332 21072
rect 14280 21029 14289 21063
rect 14289 21029 14323 21063
rect 14323 21029 14332 21063
rect 14280 21020 14332 21029
rect 10968 20884 11020 20936
rect 6460 20816 6512 20868
rect 5816 20791 5868 20800
rect 5816 20757 5825 20791
rect 5825 20757 5859 20791
rect 5859 20757 5868 20791
rect 5816 20748 5868 20757
rect 10416 20816 10468 20868
rect 10600 20816 10652 20868
rect 14096 20952 14148 21004
rect 15108 20952 15160 21004
rect 15200 20952 15252 21004
rect 12716 20884 12768 20936
rect 12808 20884 12860 20936
rect 14464 20884 14516 20936
rect 15016 20884 15068 20936
rect 18880 21020 18932 21072
rect 20812 21088 20864 21140
rect 22376 21088 22428 21140
rect 23756 21088 23808 21140
rect 24216 21131 24268 21140
rect 24216 21097 24225 21131
rect 24225 21097 24259 21131
rect 24259 21097 24268 21131
rect 24216 21088 24268 21097
rect 20260 21020 20312 21072
rect 21732 21020 21784 21072
rect 18788 20952 18840 21004
rect 20720 20952 20772 21004
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 10140 20748 10192 20800
rect 13636 20816 13688 20868
rect 13820 20816 13872 20868
rect 14280 20816 14332 20868
rect 15476 20816 15528 20868
rect 19800 20884 19852 20936
rect 22008 21020 22060 21072
rect 21916 20952 21968 21004
rect 22192 20952 22244 21004
rect 23388 20952 23440 21004
rect 23480 20952 23532 21004
rect 16764 20859 16816 20868
rect 16764 20825 16773 20859
rect 16773 20825 16807 20859
rect 16807 20825 16816 20859
rect 16764 20816 16816 20825
rect 12164 20748 12216 20800
rect 13360 20748 13412 20800
rect 14740 20748 14792 20800
rect 16672 20748 16724 20800
rect 17132 20816 17184 20868
rect 18328 20816 18380 20868
rect 19340 20816 19392 20868
rect 19616 20816 19668 20868
rect 21088 20816 21140 20868
rect 22100 20884 22152 20936
rect 23848 20884 23900 20936
rect 24308 20884 24360 20936
rect 24492 20884 24544 20936
rect 22652 20816 22704 20868
rect 24032 20816 24084 20868
rect 16948 20748 17000 20800
rect 18052 20748 18104 20800
rect 18696 20748 18748 20800
rect 20628 20748 20680 20800
rect 23388 20748 23440 20800
rect 24400 20791 24452 20800
rect 24400 20757 24409 20791
rect 24409 20757 24443 20791
rect 24443 20757 24452 20791
rect 24400 20748 24452 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 8392 20544 8444 20596
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 7104 20451 7156 20460
rect 7104 20417 7113 20451
rect 7113 20417 7147 20451
rect 7147 20417 7156 20451
rect 7104 20408 7156 20417
rect 6920 20340 6972 20392
rect 9588 20476 9640 20528
rect 10784 20544 10836 20596
rect 12256 20544 12308 20596
rect 12808 20544 12860 20596
rect 13452 20544 13504 20596
rect 14832 20544 14884 20596
rect 15200 20544 15252 20596
rect 18512 20544 18564 20596
rect 20812 20544 20864 20596
rect 11520 20476 11572 20528
rect 14280 20476 14332 20528
rect 19616 20476 19668 20528
rect 21088 20476 21140 20528
rect 10600 20408 10652 20460
rect 10876 20408 10928 20460
rect 10968 20408 11020 20460
rect 13452 20408 13504 20460
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 15936 20408 15988 20460
rect 18512 20408 18564 20460
rect 18788 20408 18840 20460
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 23296 20544 23348 20596
rect 23204 20519 23256 20528
rect 23204 20485 23213 20519
rect 23213 20485 23247 20519
rect 23247 20485 23256 20519
rect 23204 20476 23256 20485
rect 24308 20476 24360 20528
rect 9036 20383 9088 20392
rect 9036 20349 9045 20383
rect 9045 20349 9079 20383
rect 9079 20349 9088 20383
rect 9036 20340 9088 20349
rect 10692 20340 10744 20392
rect 3700 20272 3752 20324
rect 8944 20272 8996 20324
rect 7840 20204 7892 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 8484 20204 8536 20256
rect 10692 20204 10744 20256
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 15016 20340 15068 20392
rect 15200 20340 15252 20392
rect 16304 20340 16356 20392
rect 16488 20340 16540 20392
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 14924 20272 14976 20324
rect 15016 20204 15068 20256
rect 15108 20204 15160 20256
rect 17960 20204 18012 20256
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 20720 20340 20772 20392
rect 20536 20272 20588 20324
rect 22468 20340 22520 20392
rect 23388 20340 23440 20392
rect 24216 20340 24268 20392
rect 20076 20204 20128 20256
rect 20260 20204 20312 20256
rect 22376 20204 22428 20256
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 4804 20000 4856 20052
rect 7012 20000 7064 20052
rect 7932 20000 7984 20052
rect 10140 20000 10192 20052
rect 10784 20000 10836 20052
rect 4988 19932 5040 19984
rect 2872 19907 2924 19916
rect 2872 19873 2881 19907
rect 2881 19873 2915 19907
rect 2915 19873 2924 19907
rect 2872 19864 2924 19873
rect 5448 19864 5500 19916
rect 10600 19932 10652 19984
rect 3700 19796 3752 19848
rect 5908 19796 5960 19848
rect 9404 19864 9456 19916
rect 10876 19864 10928 19916
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 7472 19796 7524 19848
rect 7932 19839 7984 19848
rect 7932 19805 7941 19839
rect 7941 19805 7975 19839
rect 7975 19805 7984 19839
rect 7932 19796 7984 19805
rect 15016 20000 15068 20052
rect 17776 20000 17828 20052
rect 20260 20000 20312 20052
rect 13360 19975 13412 19984
rect 13360 19941 13369 19975
rect 13369 19941 13403 19975
rect 13403 19941 13412 19975
rect 13360 19932 13412 19941
rect 13728 19932 13780 19984
rect 13544 19864 13596 19916
rect 14280 19864 14332 19916
rect 14372 19864 14424 19916
rect 15660 19864 15712 19916
rect 18328 19932 18380 19984
rect 25044 20000 25096 20052
rect 22836 19975 22888 19984
rect 22836 19941 22845 19975
rect 22845 19941 22879 19975
rect 22879 19941 22888 19975
rect 22836 19932 22888 19941
rect 13636 19796 13688 19848
rect 13912 19796 13964 19848
rect 14556 19796 14608 19848
rect 17868 19796 17920 19848
rect 17960 19796 18012 19848
rect 22100 19864 22152 19916
rect 22652 19864 22704 19916
rect 25136 19907 25188 19916
rect 25136 19873 25145 19907
rect 25145 19873 25179 19907
rect 25179 19873 25188 19907
rect 25136 19864 25188 19873
rect 19800 19839 19852 19848
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 6092 19660 6144 19712
rect 7196 19660 7248 19712
rect 9772 19728 9824 19780
rect 11060 19728 11112 19780
rect 11888 19771 11940 19780
rect 11888 19737 11897 19771
rect 11897 19737 11931 19771
rect 11931 19737 11940 19771
rect 11888 19728 11940 19737
rect 13360 19728 13412 19780
rect 13452 19728 13504 19780
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 17500 19728 17552 19780
rect 17592 19728 17644 19780
rect 19708 19728 19760 19780
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 10784 19703 10836 19712
rect 10784 19669 10793 19703
rect 10793 19669 10827 19703
rect 10827 19669 10836 19703
rect 10784 19660 10836 19669
rect 12072 19660 12124 19712
rect 14372 19660 14424 19712
rect 16028 19660 16080 19712
rect 16304 19660 16356 19712
rect 17960 19660 18012 19712
rect 19432 19703 19484 19712
rect 19432 19669 19441 19703
rect 19441 19669 19475 19703
rect 19475 19669 19484 19703
rect 19432 19660 19484 19669
rect 19984 19660 20036 19712
rect 21088 19660 21140 19712
rect 24308 19796 24360 19848
rect 25320 19796 25372 19848
rect 23296 19660 23348 19712
rect 24492 19660 24544 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 3884 19456 3936 19508
rect 5448 19499 5500 19508
rect 5448 19465 5457 19499
rect 5457 19465 5491 19499
rect 5491 19465 5500 19499
rect 5448 19456 5500 19465
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 4804 19388 4856 19440
rect 4712 19320 4764 19372
rect 1676 19252 1728 19304
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 6184 19456 6236 19508
rect 7288 19456 7340 19508
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 6644 19388 6696 19440
rect 10416 19456 10468 19508
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 11888 19456 11940 19508
rect 14556 19456 14608 19508
rect 14832 19456 14884 19508
rect 6184 19184 6236 19236
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 6276 19116 6328 19168
rect 8484 19388 8536 19440
rect 11520 19388 11572 19440
rect 13268 19388 13320 19440
rect 13452 19388 13504 19440
rect 15016 19388 15068 19440
rect 15660 19388 15712 19440
rect 19432 19456 19484 19508
rect 20720 19456 20772 19508
rect 8024 19252 8076 19304
rect 10508 19320 10560 19372
rect 11704 19320 11756 19372
rect 12348 19320 12400 19372
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 16212 19320 16264 19372
rect 8484 19252 8536 19304
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 10692 19252 10744 19304
rect 15108 19252 15160 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 16028 19252 16080 19304
rect 10416 19184 10468 19236
rect 10784 19116 10836 19168
rect 11060 19184 11112 19236
rect 16580 19388 16632 19440
rect 17960 19388 18012 19440
rect 20536 19388 20588 19440
rect 22376 19499 22428 19508
rect 22376 19465 22385 19499
rect 22385 19465 22419 19499
rect 22419 19465 22428 19499
rect 22376 19456 22428 19465
rect 22560 19456 22612 19508
rect 25412 19456 25464 19508
rect 23664 19388 23716 19440
rect 24308 19388 24360 19440
rect 16488 19320 16540 19372
rect 16580 19252 16632 19304
rect 17684 19252 17736 19304
rect 17960 19252 18012 19304
rect 18512 19252 18564 19304
rect 19432 19320 19484 19372
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 20628 19320 20680 19372
rect 21824 19320 21876 19372
rect 13452 19116 13504 19168
rect 14556 19116 14608 19168
rect 15292 19116 15344 19168
rect 17040 19116 17092 19168
rect 19340 19184 19392 19236
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 22008 19252 22060 19304
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 25228 19252 25280 19304
rect 19524 19116 19576 19168
rect 20904 19116 20956 19168
rect 21180 19116 21232 19168
rect 22468 19116 22520 19168
rect 24768 19116 24820 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 2136 18912 2188 18964
rect 4712 18912 4764 18964
rect 4528 18844 4580 18896
rect 5632 18844 5684 18896
rect 2228 18708 2280 18760
rect 4344 18708 4396 18760
rect 5356 18776 5408 18828
rect 8392 18844 8444 18896
rect 7840 18819 7892 18828
rect 7840 18785 7849 18819
rect 7849 18785 7883 18819
rect 7883 18785 7892 18819
rect 7840 18776 7892 18785
rect 7932 18776 7984 18828
rect 8852 18844 8904 18896
rect 15384 18912 15436 18964
rect 17224 18955 17276 18964
rect 17224 18921 17233 18955
rect 17233 18921 17267 18955
rect 17267 18921 17276 18955
rect 17224 18912 17276 18921
rect 18788 18912 18840 18964
rect 19708 18912 19760 18964
rect 18420 18844 18472 18896
rect 18880 18844 18932 18896
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 8760 18708 8812 18760
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 10508 18708 10560 18760
rect 11152 18776 11204 18828
rect 11980 18776 12032 18828
rect 12348 18776 12400 18828
rect 12532 18776 12584 18828
rect 13452 18776 13504 18828
rect 14096 18776 14148 18828
rect 14924 18819 14976 18828
rect 14924 18785 14933 18819
rect 14933 18785 14967 18819
rect 14967 18785 14976 18819
rect 14924 18776 14976 18785
rect 11612 18708 11664 18760
rect 14280 18708 14332 18760
rect 16488 18776 16540 18828
rect 18328 18819 18380 18828
rect 18328 18785 18337 18819
rect 18337 18785 18371 18819
rect 18371 18785 18380 18819
rect 18328 18776 18380 18785
rect 19248 18776 19300 18828
rect 22836 18776 22888 18828
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 19892 18708 19944 18760
rect 22560 18708 22612 18760
rect 4068 18572 4120 18624
rect 8208 18640 8260 18692
rect 9404 18683 9456 18692
rect 9404 18649 9413 18683
rect 9413 18649 9447 18683
rect 9447 18649 9456 18683
rect 9404 18640 9456 18649
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 7288 18572 7340 18624
rect 9128 18572 9180 18624
rect 9496 18572 9548 18624
rect 9588 18572 9640 18624
rect 9680 18572 9732 18624
rect 11244 18640 11296 18692
rect 11520 18640 11572 18692
rect 12256 18640 12308 18692
rect 12716 18640 12768 18692
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 14556 18572 14608 18624
rect 14740 18615 14792 18624
rect 14740 18581 14749 18615
rect 14749 18581 14783 18615
rect 14783 18581 14792 18615
rect 14740 18572 14792 18581
rect 16028 18640 16080 18692
rect 15844 18572 15896 18624
rect 16212 18640 16264 18692
rect 17960 18640 18012 18692
rect 21088 18640 21140 18692
rect 24860 18844 24912 18896
rect 23848 18819 23900 18828
rect 23848 18785 23857 18819
rect 23857 18785 23891 18819
rect 23891 18785 23900 18819
rect 23848 18776 23900 18785
rect 24032 18819 24084 18828
rect 24032 18785 24041 18819
rect 24041 18785 24075 18819
rect 24075 18785 24084 18819
rect 24032 18776 24084 18785
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 24768 18708 24820 18760
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 20168 18572 20220 18624
rect 22284 18572 22336 18624
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 22928 18615 22980 18624
rect 22928 18581 22937 18615
rect 22937 18581 22971 18615
rect 22971 18581 22980 18615
rect 25320 18640 25372 18692
rect 22928 18572 22980 18581
rect 24124 18572 24176 18624
rect 25044 18615 25096 18624
rect 25044 18581 25053 18615
rect 25053 18581 25087 18615
rect 25087 18581 25096 18615
rect 25044 18572 25096 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 6828 18368 6880 18420
rect 7380 18368 7432 18420
rect 9036 18368 9088 18420
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 3332 18232 3384 18284
rect 4436 18232 4488 18284
rect 4896 18232 4948 18284
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 5264 18232 5316 18284
rect 7196 18232 7248 18284
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 8852 18300 8904 18352
rect 11152 18343 11204 18352
rect 11152 18309 11161 18343
rect 11161 18309 11195 18343
rect 11195 18309 11204 18343
rect 11152 18300 11204 18309
rect 11612 18300 11664 18352
rect 12256 18300 12308 18352
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 17316 18368 17368 18420
rect 18420 18368 18472 18420
rect 19248 18368 19300 18420
rect 20904 18368 20956 18420
rect 8668 18232 8720 18284
rect 9588 18232 9640 18284
rect 9956 18232 10008 18284
rect 11428 18232 11480 18284
rect 4620 18164 4672 18216
rect 4712 18096 4764 18148
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8392 18164 8444 18216
rect 10784 18164 10836 18216
rect 12532 18232 12584 18284
rect 18512 18300 18564 18352
rect 22744 18368 22796 18420
rect 24952 18411 25004 18420
rect 24952 18377 24961 18411
rect 24961 18377 24995 18411
rect 24995 18377 25004 18411
rect 24952 18368 25004 18377
rect 22928 18300 22980 18352
rect 15016 18232 15068 18284
rect 15568 18275 15620 18284
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 16304 18232 16356 18284
rect 17132 18232 17184 18284
rect 19892 18232 19944 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 25044 18300 25096 18352
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 14740 18164 14792 18216
rect 15660 18207 15712 18216
rect 15660 18173 15669 18207
rect 15669 18173 15703 18207
rect 15703 18173 15712 18207
rect 15660 18164 15712 18173
rect 15844 18207 15896 18216
rect 15844 18173 15853 18207
rect 15853 18173 15887 18207
rect 15887 18173 15896 18207
rect 15844 18164 15896 18173
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 20352 18164 20404 18216
rect 24768 18232 24820 18284
rect 21088 18207 21140 18216
rect 21088 18173 21097 18207
rect 21097 18173 21131 18207
rect 21131 18173 21140 18207
rect 21088 18164 21140 18173
rect 22836 18164 22888 18216
rect 5172 18139 5224 18148
rect 5172 18105 5181 18139
rect 5181 18105 5215 18139
rect 5215 18105 5224 18139
rect 5172 18096 5224 18105
rect 5724 18096 5776 18148
rect 6644 18096 6696 18148
rect 11060 18096 11112 18148
rect 12532 18096 12584 18148
rect 17224 18096 17276 18148
rect 5356 18028 5408 18080
rect 6920 18028 6972 18080
rect 9404 18028 9456 18080
rect 10600 18028 10652 18080
rect 12072 18028 12124 18080
rect 15568 18028 15620 18080
rect 16212 18028 16264 18080
rect 20628 18028 20680 18080
rect 22100 18028 22152 18080
rect 23388 18028 23440 18080
rect 23572 18028 23624 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 2044 17824 2096 17876
rect 5080 17824 5132 17876
rect 5540 17824 5592 17876
rect 7656 17824 7708 17876
rect 15844 17824 15896 17876
rect 16580 17867 16632 17876
rect 16580 17833 16589 17867
rect 16589 17833 16623 17867
rect 16623 17833 16632 17867
rect 16580 17824 16632 17833
rect 18696 17824 18748 17876
rect 21364 17824 21416 17876
rect 7104 17799 7156 17808
rect 7104 17765 7113 17799
rect 7113 17765 7147 17799
rect 7147 17765 7156 17799
rect 7104 17756 7156 17765
rect 6000 17688 6052 17740
rect 11520 17799 11572 17808
rect 11520 17765 11529 17799
rect 11529 17765 11563 17799
rect 11563 17765 11572 17799
rect 11520 17756 11572 17765
rect 13728 17799 13780 17808
rect 13728 17765 13737 17799
rect 13737 17765 13771 17799
rect 13771 17765 13780 17799
rect 13728 17756 13780 17765
rect 3792 17620 3844 17672
rect 5080 17620 5132 17672
rect 5816 17620 5868 17672
rect 3700 17552 3752 17604
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 4528 17527 4580 17536
rect 4528 17493 4537 17527
rect 4537 17493 4571 17527
rect 4571 17493 4580 17527
rect 4528 17484 4580 17493
rect 7748 17620 7800 17672
rect 9220 17620 9272 17672
rect 9680 17620 9732 17672
rect 11152 17620 11204 17672
rect 8760 17552 8812 17604
rect 9864 17484 9916 17536
rect 10968 17484 11020 17536
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12624 17688 12676 17740
rect 13452 17688 13504 17740
rect 14280 17688 14332 17740
rect 17408 17756 17460 17808
rect 21916 17824 21968 17876
rect 23388 17824 23440 17876
rect 16580 17688 16632 17740
rect 16488 17620 16540 17672
rect 19248 17620 19300 17672
rect 19616 17688 19668 17740
rect 22100 17688 22152 17740
rect 23480 17688 23532 17740
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 12716 17552 12768 17604
rect 13912 17552 13964 17604
rect 15108 17595 15160 17604
rect 15108 17561 15117 17595
rect 15117 17561 15151 17595
rect 15151 17561 15160 17595
rect 15108 17552 15160 17561
rect 15200 17552 15252 17604
rect 15568 17552 15620 17604
rect 17040 17527 17092 17536
rect 17040 17493 17049 17527
rect 17049 17493 17083 17527
rect 17083 17493 17092 17527
rect 17040 17484 17092 17493
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 17868 17484 17920 17536
rect 19708 17484 19760 17536
rect 19800 17527 19852 17536
rect 19800 17493 19809 17527
rect 19809 17493 19843 17527
rect 19843 17493 19852 17527
rect 19800 17484 19852 17493
rect 20812 17595 20864 17604
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 20904 17552 20956 17604
rect 24584 17620 24636 17672
rect 23388 17552 23440 17604
rect 22192 17484 22244 17536
rect 22744 17527 22796 17536
rect 22744 17493 22753 17527
rect 22753 17493 22787 17527
rect 22787 17493 22796 17527
rect 22744 17484 22796 17493
rect 24308 17484 24360 17536
rect 24952 17595 25004 17604
rect 24952 17561 24961 17595
rect 24961 17561 24995 17595
rect 24995 17561 25004 17595
rect 24952 17552 25004 17561
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 6736 17280 6788 17332
rect 8576 17280 8628 17332
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 9772 17280 9824 17332
rect 9864 17280 9916 17332
rect 10416 17280 10468 17332
rect 10508 17280 10560 17332
rect 3976 17144 4028 17196
rect 6092 17187 6144 17196
rect 6092 17153 6101 17187
rect 6101 17153 6135 17187
rect 6135 17153 6144 17187
rect 6092 17144 6144 17153
rect 6368 17144 6420 17196
rect 7564 17144 7616 17196
rect 7840 17144 7892 17196
rect 8852 17187 8904 17196
rect 8852 17153 8861 17187
rect 8861 17153 8895 17187
rect 8895 17153 8904 17187
rect 8852 17144 8904 17153
rect 9680 17212 9732 17264
rect 10968 17280 11020 17332
rect 11152 17212 11204 17264
rect 11060 17144 11112 17196
rect 12348 17144 12400 17196
rect 12716 17144 12768 17196
rect 17040 17280 17092 17332
rect 17224 17323 17276 17332
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 17592 17280 17644 17332
rect 19340 17280 19392 17332
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 20812 17280 20864 17332
rect 22284 17280 22336 17332
rect 22376 17280 22428 17332
rect 23296 17280 23348 17332
rect 23848 17323 23900 17332
rect 23848 17289 23857 17323
rect 23857 17289 23891 17323
rect 23891 17289 23900 17323
rect 23848 17280 23900 17289
rect 16672 17212 16724 17264
rect 17408 17212 17460 17264
rect 17776 17212 17828 17264
rect 20352 17212 20404 17264
rect 20996 17212 21048 17264
rect 6552 17076 6604 17128
rect 6828 17008 6880 17060
rect 4988 16940 5040 16992
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 10876 17076 10928 17128
rect 11980 17076 12032 17128
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 14740 17144 14792 17196
rect 15292 17144 15344 17196
rect 15844 17144 15896 17196
rect 17868 17144 17920 17196
rect 18420 17187 18472 17196
rect 18420 17153 18429 17187
rect 18429 17153 18463 17187
rect 18463 17153 18472 17187
rect 18420 17144 18472 17153
rect 20168 17144 20220 17196
rect 21456 17187 21508 17196
rect 21456 17153 21465 17187
rect 21465 17153 21499 17187
rect 21499 17153 21508 17187
rect 21456 17144 21508 17153
rect 10600 17008 10652 17060
rect 16212 17119 16264 17128
rect 16212 17085 16221 17119
rect 16221 17085 16255 17119
rect 16255 17085 16264 17119
rect 16212 17076 16264 17085
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 20996 17076 21048 17128
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 23480 17144 23532 17196
rect 13360 16983 13412 16992
rect 13360 16949 13369 16983
rect 13369 16949 13403 16983
rect 13403 16949 13412 16983
rect 13360 16940 13412 16949
rect 16580 16940 16632 16992
rect 17040 16940 17092 16992
rect 21916 17008 21968 17060
rect 21180 16940 21232 16992
rect 21732 16940 21784 16992
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 25412 17212 25464 17264
rect 23940 17008 23992 17060
rect 23756 16940 23808 16992
rect 25412 17008 25464 17060
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 4896 16779 4948 16788
rect 4896 16745 4905 16779
rect 4905 16745 4939 16779
rect 4939 16745 4948 16779
rect 4896 16736 4948 16745
rect 4988 16736 5040 16788
rect 9956 16736 10008 16788
rect 10232 16736 10284 16788
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 6736 16711 6788 16720
rect 6736 16677 6745 16711
rect 6745 16677 6779 16711
rect 6779 16677 6788 16711
rect 6736 16668 6788 16677
rect 7472 16668 7524 16720
rect 9220 16668 9272 16720
rect 8944 16532 8996 16584
rect 14096 16668 14148 16720
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 17592 16736 17644 16788
rect 19432 16736 19484 16788
rect 10968 16600 11020 16652
rect 13728 16600 13780 16652
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 17040 16668 17092 16720
rect 20996 16736 21048 16788
rect 21364 16668 21416 16720
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 16856 16600 16908 16652
rect 19340 16600 19392 16652
rect 22100 16600 22152 16652
rect 23572 16600 23624 16652
rect 24584 16600 24636 16652
rect 11060 16532 11112 16584
rect 11704 16532 11756 16584
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 5172 16464 5224 16516
rect 12532 16464 12584 16516
rect 12716 16464 12768 16516
rect 15292 16464 15344 16516
rect 17868 16464 17920 16516
rect 18696 16464 18748 16516
rect 20168 16464 20220 16516
rect 23572 16464 23624 16516
rect 24676 16507 24728 16516
rect 24676 16473 24685 16507
rect 24685 16473 24719 16507
rect 24719 16473 24728 16507
rect 24676 16464 24728 16473
rect 6092 16439 6144 16448
rect 6092 16405 6101 16439
rect 6101 16405 6135 16439
rect 6135 16405 6144 16439
rect 6092 16396 6144 16405
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 9956 16396 10008 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 12072 16396 12124 16448
rect 17316 16396 17368 16448
rect 21272 16396 21324 16448
rect 21456 16396 21508 16448
rect 22008 16396 22060 16448
rect 23940 16396 23992 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 9128 16235 9180 16244
rect 9128 16201 9137 16235
rect 9137 16201 9171 16235
rect 9171 16201 9180 16235
rect 9128 16192 9180 16201
rect 9220 16192 9272 16244
rect 10968 16235 11020 16244
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 11520 16192 11572 16244
rect 16212 16192 16264 16244
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 18972 16192 19024 16244
rect 19248 16192 19300 16244
rect 5172 16099 5224 16108
rect 5172 16065 5181 16099
rect 5181 16065 5215 16099
rect 5215 16065 5224 16099
rect 5172 16056 5224 16065
rect 8576 16056 8628 16108
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 4252 15988 4304 16040
rect 11060 16124 11112 16176
rect 12072 16124 12124 16176
rect 12256 16124 12308 16176
rect 12440 16124 12492 16176
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 21824 16192 21876 16244
rect 22008 16192 22060 16244
rect 24400 16192 24452 16244
rect 20444 16124 20496 16176
rect 10232 16056 10284 16108
rect 14096 16056 14148 16108
rect 15844 16056 15896 16108
rect 17132 16056 17184 16108
rect 17960 16056 18012 16108
rect 18696 16056 18748 16108
rect 10140 15988 10192 16040
rect 10508 15988 10560 16040
rect 10600 15988 10652 16040
rect 6092 15920 6144 15972
rect 10968 15988 11020 16040
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12072 15988 12124 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 15660 15988 15712 16040
rect 7012 15852 7064 15904
rect 10600 15852 10652 15904
rect 15568 15963 15620 15972
rect 15568 15929 15577 15963
rect 15577 15929 15611 15963
rect 15611 15929 15620 15963
rect 15568 15920 15620 15929
rect 13820 15852 13872 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 14648 15852 14700 15904
rect 16764 15988 16816 16040
rect 20996 16056 21048 16108
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 21640 16056 21692 16108
rect 24216 16056 24268 16108
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 22284 15988 22336 16040
rect 23940 16031 23992 16040
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 17040 15920 17092 15972
rect 18972 15852 19024 15904
rect 21640 15852 21692 15904
rect 22376 15852 22428 15904
rect 25228 15920 25280 15972
rect 25136 15852 25188 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 8484 15648 8536 15700
rect 13912 15648 13964 15700
rect 15108 15648 15160 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 22468 15648 22520 15700
rect 10232 15580 10284 15632
rect 12072 15580 12124 15632
rect 19984 15580 20036 15632
rect 11520 15512 11572 15564
rect 13728 15512 13780 15564
rect 16488 15512 16540 15564
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 20260 15512 20312 15564
rect 22560 15580 22612 15632
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 10324 15444 10376 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 20536 15444 20588 15496
rect 22284 15444 22336 15496
rect 23664 15444 23716 15496
rect 12348 15376 12400 15428
rect 13360 15376 13412 15428
rect 15292 15376 15344 15428
rect 17316 15376 17368 15428
rect 17776 15376 17828 15428
rect 19800 15376 19852 15428
rect 21180 15376 21232 15428
rect 11796 15308 11848 15360
rect 11980 15308 12032 15360
rect 16580 15308 16632 15360
rect 17224 15308 17276 15360
rect 19892 15308 19944 15360
rect 21732 15308 21784 15360
rect 22836 15351 22888 15360
rect 22836 15317 22845 15351
rect 22845 15317 22879 15351
rect 22879 15317 22888 15351
rect 22836 15308 22888 15317
rect 23296 15308 23348 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 11244 15104 11296 15156
rect 12072 15104 12124 15156
rect 15384 15104 15436 15156
rect 16764 15104 16816 15156
rect 16856 15104 16908 15156
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 11888 15036 11940 15088
rect 12440 15036 12492 15088
rect 13912 15036 13964 15088
rect 17224 15036 17276 15088
rect 17776 15036 17828 15088
rect 21364 15104 21416 15156
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 25044 15104 25096 15156
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 20996 15036 21048 15088
rect 21272 15036 21324 15088
rect 22652 15036 22704 15088
rect 23664 15036 23716 15088
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 10692 14900 10744 14952
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 12440 14900 12492 14952
rect 14648 14900 14700 14952
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 15476 14900 15528 14952
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 25320 15011 25372 15020
rect 25320 14977 25329 15011
rect 25329 14977 25363 15011
rect 25363 14977 25372 15011
rect 25320 14968 25372 14977
rect 18788 14900 18840 14952
rect 19708 14943 19760 14952
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 21916 14900 21968 14952
rect 23940 14900 23992 14952
rect 16672 14832 16724 14884
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 18880 14832 18932 14884
rect 22468 14832 22520 14884
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 10600 14560 10652 14612
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 12808 14560 12860 14612
rect 13360 14560 13412 14612
rect 13820 14560 13872 14612
rect 15016 14560 15068 14612
rect 15660 14560 15712 14612
rect 23388 14560 23440 14612
rect 14004 14492 14056 14544
rect 16488 14492 16540 14544
rect 18328 14492 18380 14544
rect 18788 14492 18840 14544
rect 21180 14492 21232 14544
rect 11980 14424 12032 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 18604 14424 18656 14476
rect 12348 14288 12400 14340
rect 14556 14331 14608 14340
rect 14556 14297 14565 14331
rect 14565 14297 14599 14331
rect 14599 14297 14608 14331
rect 14556 14288 14608 14297
rect 15292 14288 15344 14340
rect 12716 14220 12768 14272
rect 14832 14220 14884 14272
rect 19892 14356 19944 14408
rect 24032 14424 24084 14476
rect 25044 14356 25096 14408
rect 16672 14288 16724 14340
rect 17040 14220 17092 14272
rect 17316 14288 17368 14340
rect 18512 14288 18564 14340
rect 20904 14288 20956 14340
rect 23572 14288 23624 14340
rect 24492 14288 24544 14340
rect 25596 14288 25648 14340
rect 19064 14220 19116 14272
rect 19524 14220 19576 14272
rect 21916 14220 21968 14272
rect 23848 14220 23900 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 13452 14016 13504 14068
rect 14188 14016 14240 14068
rect 14556 14016 14608 14068
rect 15844 14016 15896 14068
rect 17224 14016 17276 14068
rect 17684 14016 17736 14068
rect 19432 14016 19484 14068
rect 20996 14016 21048 14068
rect 23480 14016 23532 14068
rect 23572 14016 23624 14068
rect 12808 13880 12860 13932
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 14280 13948 14332 14000
rect 15292 13948 15344 14000
rect 17592 13948 17644 14000
rect 18328 13948 18380 14000
rect 18512 13948 18564 14000
rect 19064 13948 19116 14000
rect 20904 13948 20956 14000
rect 16488 13880 16540 13932
rect 17316 13880 17368 13932
rect 18420 13880 18472 13932
rect 20720 13880 20772 13932
rect 13912 13812 13964 13864
rect 14372 13812 14424 13864
rect 17592 13812 17644 13864
rect 16028 13744 16080 13796
rect 17776 13812 17828 13864
rect 23664 13880 23716 13932
rect 15568 13676 15620 13728
rect 19708 13744 19760 13796
rect 21916 13812 21968 13864
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 24492 13855 24544 13864
rect 24492 13821 24501 13855
rect 24501 13821 24535 13855
rect 24535 13821 24544 13855
rect 24492 13812 24544 13821
rect 21456 13744 21508 13796
rect 21548 13744 21600 13796
rect 22192 13744 22244 13796
rect 20168 13676 20220 13728
rect 20352 13676 20404 13728
rect 21364 13676 21416 13728
rect 21732 13676 21784 13728
rect 24676 13676 24728 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 13176 13472 13228 13524
rect 17408 13472 17460 13524
rect 18880 13515 18932 13524
rect 18880 13481 18889 13515
rect 18889 13481 18923 13515
rect 18923 13481 18932 13515
rect 18880 13472 18932 13481
rect 15568 13404 15620 13456
rect 20076 13472 20128 13524
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 16948 13336 17000 13388
rect 19156 13336 19208 13388
rect 19432 13336 19484 13388
rect 20352 13336 20404 13388
rect 20536 13336 20588 13388
rect 24860 13336 24912 13388
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 9588 13311 9640 13320
rect 9588 13277 9597 13311
rect 9597 13277 9631 13311
rect 9631 13277 9640 13311
rect 9588 13268 9640 13277
rect 10140 13132 10192 13184
rect 10692 13132 10744 13184
rect 21916 13311 21968 13320
rect 21916 13277 21925 13311
rect 21925 13277 21959 13311
rect 21959 13277 21968 13311
rect 21916 13268 21968 13277
rect 13728 13200 13780 13252
rect 14648 13200 14700 13252
rect 12440 13132 12492 13184
rect 13636 13132 13688 13184
rect 15292 13132 15344 13184
rect 16488 13200 16540 13252
rect 18972 13200 19024 13252
rect 19156 13200 19208 13252
rect 21272 13200 21324 13252
rect 21364 13200 21416 13252
rect 16304 13132 16356 13184
rect 21548 13132 21600 13184
rect 22192 13243 22244 13252
rect 22192 13209 22201 13243
rect 22201 13209 22235 13243
rect 22235 13209 22244 13243
rect 22192 13200 22244 13209
rect 22652 13200 22704 13252
rect 23572 13200 23624 13252
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 14188 12928 14240 12980
rect 14648 12971 14700 12980
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 13176 12903 13228 12912
rect 13176 12869 13185 12903
rect 13185 12869 13219 12903
rect 13219 12869 13228 12903
rect 13176 12860 13228 12869
rect 13636 12860 13688 12912
rect 18328 12860 18380 12912
rect 17868 12792 17920 12844
rect 19432 12928 19484 12980
rect 19800 12928 19852 12980
rect 22192 12928 22244 12980
rect 25136 12928 25188 12980
rect 18788 12903 18840 12912
rect 18788 12869 18797 12903
rect 18797 12869 18831 12903
rect 18831 12869 18840 12903
rect 18788 12860 18840 12869
rect 20076 12860 20128 12912
rect 21272 12860 21324 12912
rect 22928 12860 22980 12912
rect 18236 12724 18288 12776
rect 25044 12835 25096 12844
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 20168 12656 20220 12708
rect 20812 12656 20864 12708
rect 23480 12724 23532 12776
rect 23940 12656 23992 12708
rect 24676 12656 24728 12708
rect 17040 12588 17092 12640
rect 18604 12588 18656 12640
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 20444 12588 20496 12640
rect 23020 12588 23072 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 16672 12384 16724 12436
rect 4160 12248 4212 12300
rect 17040 12248 17092 12300
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 18420 12384 18472 12436
rect 19524 12384 19576 12436
rect 19708 12427 19760 12436
rect 19708 12393 19738 12427
rect 19738 12393 19760 12427
rect 19708 12384 19760 12393
rect 21088 12384 21140 12436
rect 21364 12384 21416 12436
rect 21732 12384 21784 12436
rect 17224 12316 17276 12368
rect 24216 12384 24268 12436
rect 24676 12316 24728 12368
rect 20720 12248 20772 12300
rect 18328 12180 18380 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 16028 12155 16080 12164
rect 16028 12121 16037 12155
rect 16037 12121 16071 12155
rect 16071 12121 16080 12155
rect 16028 12112 16080 12121
rect 19340 12112 19392 12164
rect 20168 12112 20220 12164
rect 21088 12248 21140 12300
rect 24032 12248 24084 12300
rect 21180 12180 21232 12232
rect 22008 12180 22060 12232
rect 22652 12112 22704 12164
rect 19616 12044 19668 12096
rect 21088 12044 21140 12096
rect 21456 12044 21508 12096
rect 21640 12087 21692 12096
rect 21640 12053 21649 12087
rect 21649 12053 21683 12087
rect 21683 12053 21692 12087
rect 21640 12044 21692 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 14464 11883 14516 11892
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 15844 11883 15896 11892
rect 15844 11849 15853 11883
rect 15853 11849 15887 11883
rect 15887 11849 15896 11883
rect 15844 11840 15896 11849
rect 15936 11840 15988 11892
rect 19248 11840 19300 11892
rect 16580 11772 16632 11824
rect 15844 11704 15896 11756
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 17040 11772 17092 11824
rect 17224 11772 17276 11824
rect 18144 11772 18196 11824
rect 21180 11840 21232 11892
rect 19616 11815 19668 11824
rect 19616 11781 19625 11815
rect 19625 11781 19659 11815
rect 19659 11781 19668 11815
rect 19616 11772 19668 11781
rect 20076 11772 20128 11824
rect 24860 11772 24912 11824
rect 21640 11704 21692 11756
rect 14556 11636 14608 11688
rect 20076 11636 20128 11688
rect 20260 11636 20312 11688
rect 21548 11636 21600 11688
rect 21916 11636 21968 11688
rect 23480 11704 23532 11756
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 14280 11568 14332 11620
rect 16856 11568 16908 11620
rect 17684 11500 17736 11552
rect 20628 11500 20680 11552
rect 21088 11500 21140 11552
rect 24584 11500 24636 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 6552 11296 6604 11348
rect 16396 11296 16448 11348
rect 19708 11228 19760 11280
rect 19432 11160 19484 11212
rect 16948 11092 17000 11144
rect 20996 11296 21048 11348
rect 22008 11296 22060 11348
rect 23940 11296 23992 11348
rect 24584 11339 24636 11348
rect 24584 11305 24593 11339
rect 24593 11305 24627 11339
rect 24627 11305 24636 11339
rect 24584 11296 24636 11305
rect 24032 11228 24084 11280
rect 20076 11160 20128 11212
rect 20168 11160 20220 11212
rect 17684 11024 17736 11076
rect 18144 11024 18196 11076
rect 20628 11024 20680 11076
rect 21272 11092 21324 11144
rect 21824 11092 21876 11144
rect 24952 11160 25004 11212
rect 24400 11092 24452 11144
rect 18420 10956 18472 11008
rect 18880 10956 18932 11008
rect 21732 11024 21784 11076
rect 23296 11024 23348 11076
rect 22008 10956 22060 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 16764 10752 16816 10804
rect 18512 10752 18564 10804
rect 18880 10752 18932 10804
rect 17592 10684 17644 10736
rect 10232 10616 10284 10668
rect 17316 10616 17368 10668
rect 17776 10616 17828 10668
rect 17960 10684 18012 10736
rect 20812 10684 20864 10736
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 19248 10616 19300 10668
rect 19800 10616 19852 10668
rect 20536 10616 20588 10668
rect 20904 10659 20956 10668
rect 20904 10625 20913 10659
rect 20913 10625 20947 10659
rect 20947 10625 20956 10659
rect 20904 10616 20956 10625
rect 24860 10684 24912 10736
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 20168 10548 20220 10600
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 19984 10480 20036 10532
rect 25136 10480 25188 10532
rect 19432 10455 19484 10464
rect 19432 10421 19441 10455
rect 19441 10421 19475 10455
rect 19475 10421 19484 10455
rect 19432 10412 19484 10421
rect 20168 10412 20220 10464
rect 21364 10412 21416 10464
rect 22284 10412 22336 10464
rect 22744 10412 22796 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 17500 10208 17552 10260
rect 19524 10208 19576 10260
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 20720 10140 20772 10192
rect 20260 10072 20312 10124
rect 20076 10004 20128 10056
rect 21180 10072 21232 10124
rect 21548 10115 21600 10124
rect 21548 10081 21557 10115
rect 21557 10081 21591 10115
rect 21591 10081 21600 10115
rect 21548 10072 21600 10081
rect 22192 10072 22244 10124
rect 20536 10004 20588 10056
rect 20720 9936 20772 9988
rect 22652 10004 22704 10056
rect 24124 10004 24176 10056
rect 21824 9936 21876 9988
rect 23940 9936 23992 9988
rect 23020 9911 23072 9920
rect 23020 9877 23029 9911
rect 23029 9877 23063 9911
rect 23063 9877 23072 9911
rect 25044 10004 25096 10056
rect 23020 9868 23072 9877
rect 25136 9868 25188 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 20076 9664 20128 9716
rect 20536 9664 20588 9716
rect 17408 9596 17460 9648
rect 20720 9664 20772 9716
rect 21824 9664 21876 9716
rect 23020 9664 23072 9716
rect 18696 9528 18748 9580
rect 18972 9528 19024 9580
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 16120 9392 16172 9444
rect 22376 9460 22428 9512
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 18696 9367 18748 9376
rect 18696 9333 18705 9367
rect 18705 9333 18739 9367
rect 18739 9333 18748 9367
rect 18696 9324 18748 9333
rect 20260 9324 20312 9376
rect 24308 9392 24360 9444
rect 23388 9324 23440 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 14372 9120 14424 9172
rect 19524 9120 19576 9172
rect 26056 9120 26108 9172
rect 16856 9052 16908 9104
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 18696 8984 18748 9036
rect 20812 8916 20864 8968
rect 25688 9052 25740 9104
rect 24952 8984 25004 9036
rect 6828 8848 6880 8900
rect 12348 8848 12400 8900
rect 22560 8916 22612 8968
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 24400 8848 24452 8900
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 25136 8848 25188 8900
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 14740 8576 14792 8628
rect 23480 8576 23532 8628
rect 20352 8508 20404 8560
rect 20444 8440 20496 8492
rect 20720 8508 20772 8560
rect 21732 8440 21784 8492
rect 24860 8508 24912 8560
rect 25228 8440 25280 8492
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 24032 8304 24084 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 22652 8032 22704 8084
rect 24400 8032 24452 8084
rect 21916 7964 21968 8016
rect 23572 7964 23624 8016
rect 21640 7896 21692 7948
rect 19432 7828 19484 7880
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 24952 7896 25004 7948
rect 24860 7760 24912 7812
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 25412 7488 25464 7540
rect 24860 7420 24912 7472
rect 23388 7352 23440 7404
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 25044 7216 25096 7268
rect 22744 7148 22796 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 21364 6740 21416 6792
rect 22284 6740 22336 6792
rect 24860 6808 24912 6860
rect 24308 6740 24360 6792
rect 11612 6672 11664 6724
rect 25044 6672 25096 6724
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 25136 6400 25188 6452
rect 24860 6332 24912 6384
rect 24492 6264 24544 6316
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 23296 5788 23348 5840
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 24124 5652 24176 5704
rect 24952 5584 25004 5636
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 20812 5244 20864 5296
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 24860 5244 24912 5296
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 22468 4564 22520 4616
rect 24032 4564 24084 4616
rect 24952 4496 25004 4548
rect 24676 4471 24728 4480
rect 24676 4437 24685 4471
rect 24685 4437 24719 4471
rect 24719 4437 24728 4471
rect 24676 4428 24728 4437
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 21180 4088 21232 4140
rect 17132 4020 17184 4072
rect 20168 4020 20220 4072
rect 22192 4020 22244 4072
rect 22836 4088 22888 4140
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 25044 3884 25096 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 22744 3544 22796 3596
rect 20628 3476 20680 3528
rect 24676 3476 24728 3528
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 24952 3408 25004 3460
rect 22284 3340 22336 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 24860 3068 24912 3120
rect 25136 3111 25188 3120
rect 25136 3077 25145 3111
rect 25145 3077 25179 3111
rect 25179 3077 25188 3111
rect 25136 3068 25188 3077
rect 18788 3000 18840 3052
rect 19340 3000 19392 3052
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 23848 3000 23900 3052
rect 19524 2932 19576 2984
rect 25044 2932 25096 2984
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 6828 2635 6880 2644
rect 6828 2601 6837 2635
rect 6837 2601 6871 2635
rect 6871 2601 6880 2635
rect 6828 2592 6880 2601
rect 23388 2456 23440 2508
rect 6736 2388 6788 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 19524 2320 19576 2372
rect 22100 2320 22152 2372
rect 23296 2388 23348 2440
rect 24952 2320 25004 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1674 26200 1730 27000
rect 2042 26200 2098 27000
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 2410 26330 2466 27000
rect 2778 26466 2834 27000
rect 2778 26450 3096 26466
rect 2778 26444 3108 26450
rect 2778 26438 3056 26444
rect 938 23760 994 23769
rect 938 23695 940 23704
rect 992 23695 994 23704
rect 940 23666 992 23672
rect 938 22672 994 22681
rect 938 22607 940 22616
rect 992 22607 994 22616
rect 940 22578 992 22584
rect 1688 19310 1716 26200
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 19378 1992 22918
rect 2056 22166 2084 26200
rect 2134 24984 2190 24993
rect 2134 24919 2190 24928
rect 2044 22160 2096 22166
rect 2044 22102 2096 22108
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 2056 18290 2084 21082
rect 2148 18970 2176 24919
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2240 18766 2268 26318
rect 2410 26302 2728 26330
rect 2410 26200 2466 26302
rect 2700 21570 2728 26302
rect 2778 26200 2834 26438
rect 3056 26386 3108 26392
rect 3146 26330 3202 27000
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 2884 26302 3202 26330
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 21690 2820 25871
rect 2884 22098 2912 26302
rect 3146 26200 3202 26302
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2700 21542 2820 21570
rect 2792 21078 2820 21542
rect 2976 21332 3004 22102
rect 2884 21304 3004 21332
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2884 19922 2912 21304
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 3344 20398 3372 26386
rect 3514 26200 3570 27000
rect 3882 26330 3938 27000
rect 3882 26302 4108 26330
rect 3882 26200 3938 26302
rect 3422 24848 3478 24857
rect 3422 24783 3478 24792
rect 3436 22030 3464 24783
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3528 21486 3556 26200
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3608 23112 3660 23118
rect 3608 23054 3660 23060
rect 3620 22166 3648 23054
rect 3608 22160 3660 22166
rect 3608 22102 3660 22108
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3712 20330 3740 24006
rect 3790 23080 3846 23089
rect 3790 23015 3846 23024
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3330 19000 3386 19009
rect 3330 18935 3386 18944
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 3344 18290 3372 18935
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 2056 17882 2084 18226
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 3238 17640 3294 17649
rect 3712 17610 3740 19790
rect 3804 17678 3832 23015
rect 3896 19514 3924 24142
rect 4080 22094 4108 26302
rect 4250 26200 4306 27000
rect 4618 26200 4674 27000
rect 4986 26200 5042 27000
rect 5354 26330 5410 27000
rect 5092 26302 5410 26330
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 23866 4200 24142
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4172 22982 4200 23258
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4264 22710 4292 26200
rect 4526 24304 4582 24313
rect 4526 24239 4582 24248
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4356 23118 4384 23530
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4540 22794 4568 24239
rect 4632 23186 4660 26200
rect 4896 24676 4948 24682
rect 4896 24618 4948 24624
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4816 24206 4844 24550
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4908 23730 4936 24618
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4710 23216 4766 23225
rect 4620 23180 4672 23186
rect 4710 23151 4766 23160
rect 4620 23122 4672 23128
rect 4356 22766 4568 22794
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4356 22522 4384 22766
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4264 22494 4384 22522
rect 4080 22066 4200 22094
rect 4172 21010 4200 22066
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 3974 19952 4030 19961
rect 3974 19887 4030 19896
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3238 17575 3294 17584
rect 3700 17604 3752 17610
rect 3252 17542 3280 17575
rect 3700 17546 3752 17552
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3988 17202 4016 19887
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 4080 14634 4108 18566
rect 4264 16046 4292 22494
rect 4448 22420 4476 22646
rect 4528 22636 4580 22642
rect 4528 22578 4580 22584
rect 4540 22522 4568 22578
rect 4540 22494 4660 22522
rect 4342 22400 4398 22409
rect 4448 22392 4568 22420
rect 4342 22335 4398 22344
rect 4356 18766 4384 22335
rect 4434 22264 4490 22273
rect 4434 22199 4490 22208
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4448 18290 4476 22199
rect 4540 22030 4568 22392
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 18902 4568 21830
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4632 18222 4660 22494
rect 4724 22273 4752 23151
rect 4710 22264 4766 22273
rect 4710 22199 4766 22208
rect 4804 22024 4856 22030
rect 4856 21984 4936 22012
rect 4804 21966 4856 21972
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 19378 4752 21830
rect 4802 21584 4858 21593
rect 4802 21519 4804 21528
rect 4856 21519 4858 21528
rect 4804 21490 4856 21496
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4816 19446 4844 19994
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18970 4752 19110
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4908 18290 4936 21984
rect 5000 21486 5028 26200
rect 5092 23798 5120 26302
rect 5264 26240 5316 26246
rect 5354 26200 5410 26302
rect 5446 26208 5502 26217
rect 5264 26182 5316 26188
rect 5170 24848 5226 24857
rect 5170 24783 5226 24792
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 5080 23248 5132 23254
rect 5080 23190 5132 23196
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 5000 18290 5028 19926
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4710 18184 4766 18193
rect 4710 18119 4712 18128
rect 4764 18119 4766 18128
rect 4712 18090 4764 18096
rect 5092 17882 5120 23190
rect 5184 22642 5212 24783
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5170 20360 5226 20369
rect 5170 20295 5226 20304
rect 5184 18154 5212 20295
rect 5276 18290 5304 26182
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26200 6514 27000
rect 6826 26200 6882 27000
rect 7194 26200 7250 27000
rect 7562 26200 7618 27000
rect 7930 26330 7986 27000
rect 7668 26302 7986 26330
rect 5446 26143 5502 26152
rect 5460 24290 5488 26143
rect 5368 24262 5488 24290
rect 5368 23254 5396 24262
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5460 19922 5488 24142
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 5540 22024 5592 22030
rect 5644 22001 5672 23054
rect 5736 22710 5764 26200
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 6104 22098 6132 26200
rect 6472 24274 6500 26200
rect 6552 24744 6604 24750
rect 6552 24686 6604 24692
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6564 23730 6592 24686
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6552 23520 6604 23526
rect 6748 23497 6776 23598
rect 6552 23462 6604 23468
rect 6734 23488 6790 23497
rect 6564 22681 6592 23462
rect 6840 23474 6868 26200
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7024 23526 7052 24142
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7012 23520 7064 23526
rect 6840 23446 6960 23474
rect 7012 23462 7064 23468
rect 6734 23423 6790 23432
rect 6550 22672 6606 22681
rect 6550 22607 6606 22616
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 5540 21966 5592 21972
rect 5630 21992 5686 22001
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5460 19417 5488 19450
rect 5446 19408 5502 19417
rect 5446 19343 5502 19352
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5368 18086 5396 18770
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5552 17882 5580 21966
rect 5630 21927 5686 21936
rect 6182 21448 6238 21457
rect 6182 21383 6238 21392
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5998 20904 6054 20913
rect 5630 20632 5686 20641
rect 5630 20567 5686 20576
rect 5644 19378 5672 20567
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5630 19272 5686 19281
rect 5630 19207 5686 19216
rect 5644 18902 5672 19207
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5736 18154 5764 20878
rect 5998 20839 6054 20848
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5092 17678 5120 17818
rect 5828 17678 5856 20742
rect 6012 20466 6040 20839
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5920 19360 5948 19790
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 5920 19332 6040 19360
rect 6012 17746 6040 19332
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4540 16153 4568 17478
rect 4894 17232 4950 17241
rect 6104 17202 6132 19654
rect 6196 19514 6224 21383
rect 6366 21176 6422 21185
rect 6366 21111 6422 21120
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6196 19242 6224 19450
rect 6184 19236 6236 19242
rect 6184 19178 6236 19184
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 4894 17167 4950 17176
rect 6092 17196 6144 17202
rect 4908 16794 4936 17167
rect 6092 17138 6144 17144
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16794 5028 16934
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 6288 16561 6316 19110
rect 6380 17202 6408 21111
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 20505 6500 20810
rect 6458 20496 6514 20505
rect 6458 20431 6514 20440
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6564 17134 6592 20878
rect 6656 19446 6684 22578
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6748 21622 6776 22374
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 6644 18760 6696 18766
rect 6840 18714 6868 22578
rect 6932 21078 6960 23446
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 7024 21078 7052 22442
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 7116 20466 7144 24006
rect 7208 21486 7236 26200
rect 7576 23798 7604 26200
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 19825 6960 20334
rect 7102 20224 7158 20233
rect 7102 20159 7158 20168
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6918 19816 6974 19825
rect 6918 19751 6974 19760
rect 6918 19544 6974 19553
rect 6918 19479 6974 19488
rect 6644 18702 6696 18708
rect 6656 18154 6684 18702
rect 6748 18686 6868 18714
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6748 17338 6776 18686
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6840 18329 6868 18362
rect 6826 18320 6882 18329
rect 6826 18255 6882 18264
rect 6932 18170 6960 19479
rect 6840 18142 6960 18170
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6840 17218 6868 18142
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6748 17190 6868 17218
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6274 16552 6330 16561
rect 5172 16516 5224 16522
rect 6274 16487 6330 16496
rect 5172 16458 5224 16464
rect 4526 16144 4582 16153
rect 5184 16114 5212 16458
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 4526 16079 4582 16088
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 6104 15978 6132 16390
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 4080 14606 4200 14634
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 4172 12306 4200 14606
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 6564 11354 6592 16934
rect 6748 16726 6776 17190
rect 6826 17096 6882 17105
rect 6826 17031 6828 17040
rect 6880 17031 6882 17040
rect 6828 17002 6880 17008
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6932 15473 6960 18022
rect 7024 15910 7052 19994
rect 7116 19553 7144 20159
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7102 19544 7158 19553
rect 7102 19479 7158 19488
rect 7102 18728 7158 18737
rect 7102 18663 7158 18672
rect 7116 18630 7144 18663
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7208 18290 7236 19654
rect 7300 19514 7328 23666
rect 7470 23624 7526 23633
rect 7470 23559 7526 23568
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 18290 7328 18566
rect 7392 18426 7420 23122
rect 7484 22030 7512 23559
rect 7668 23254 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26200 8722 27000
rect 9034 26330 9090 27000
rect 8772 26302 9090 26330
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7656 23248 7708 23254
rect 7656 23190 7708 23196
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7562 22536 7618 22545
rect 7562 22471 7618 22480
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7104 17808 7156 17814
rect 7102 17776 7104 17785
rect 7156 17776 7158 17785
rect 7102 17711 7158 17720
rect 7484 16726 7512 19790
rect 7576 17202 7604 22471
rect 7760 21146 7788 22578
rect 8312 22098 8340 26200
rect 8574 24712 8630 24721
rect 8574 24647 8630 24656
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7852 21049 7880 21830
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7838 21040 7894 21049
rect 7838 20975 7894 20984
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 17882 7696 20878
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8404 20602 8432 23666
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8496 22953 8524 23598
rect 8588 23338 8616 24647
rect 8680 24138 8708 26200
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8588 23310 8708 23338
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8482 22944 8538 22953
rect 8482 22879 8538 22888
rect 8588 22778 8616 23122
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7760 17678 7788 19450
rect 7852 19334 7880 20198
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7944 19854 7972 19994
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7852 19306 7972 19334
rect 7838 18864 7894 18873
rect 7944 18834 7972 19306
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 7838 18799 7840 18808
rect 7892 18799 7894 18808
rect 7932 18828 7984 18834
rect 7840 18770 7892 18776
rect 7932 18770 7984 18776
rect 8036 18612 8064 19246
rect 8404 18902 8432 20198
rect 8496 19446 8524 20198
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8208 18692 8260 18698
rect 8260 18652 8432 18680
rect 8208 18634 8260 18640
rect 7852 18584 8064 18612
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7852 17202 7880 18584
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8404 18465 8432 18652
rect 8390 18456 8446 18465
rect 8390 18391 8446 18400
rect 7932 18216 7984 18222
rect 8392 18216 8444 18222
rect 7932 18158 7984 18164
rect 8390 18184 8392 18193
rect 8444 18184 8446 18193
rect 7944 17921 7972 18158
rect 8390 18119 8446 18128
rect 8390 18048 8446 18057
rect 8390 17983 8446 17992
rect 7930 17912 7986 17921
rect 7930 17847 7986 17856
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 8404 16454 8432 17983
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 8496 15706 8524 19246
rect 8588 17338 8616 21490
rect 8680 18290 8708 23310
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 9692 26302 9826 26330
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23769 9168 24006
rect 9126 23760 9182 23769
rect 9126 23695 9182 23704
rect 8942 23488 8998 23497
rect 8942 23423 8998 23432
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8758 22264 8814 22273
rect 8758 22199 8814 22208
rect 8772 18766 8800 22199
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8864 19009 8892 21830
rect 8956 20330 8984 23423
rect 9416 23254 9444 26200
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 10138 26200 10194 27000
rect 10506 26200 10562 27000
rect 10874 26200 10930 27000
rect 11242 26330 11298 27000
rect 11072 26302 11298 26330
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 9140 22098 9168 22510
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 9140 21486 9168 22034
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9036 20392 9088 20398
rect 9140 20380 9168 21422
rect 9324 20942 9352 22374
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9218 20632 9274 20641
rect 9218 20567 9274 20576
rect 9088 20352 9168 20380
rect 9036 20334 9088 20340
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 8942 19544 8998 19553
rect 8942 19479 8998 19488
rect 8850 19000 8906 19009
rect 8850 18935 8906 18944
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8864 18358 8892 18838
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8668 18284 8720 18290
rect 8720 18244 8800 18272
rect 8668 18226 8720 18232
rect 8666 18184 8722 18193
rect 8666 18119 8722 18128
rect 8680 17338 8708 18119
rect 8772 17921 8800 18244
rect 8758 17912 8814 17921
rect 8758 17847 8814 17856
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8574 16280 8630 16289
rect 8574 16215 8630 16224
rect 8588 16114 8616 16215
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 6918 15464 6974 15473
rect 6918 15399 6974 15408
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8772 14385 8800 17546
rect 8850 17232 8906 17241
rect 8850 17167 8852 17176
rect 8904 17167 8906 17176
rect 8852 17138 8904 17144
rect 8956 16590 8984 19479
rect 9140 19310 9168 20352
rect 9232 20233 9260 20567
rect 9218 20224 9274 20233
rect 9218 20159 9274 20168
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 19009 9168 19246
rect 9218 19136 9274 19145
rect 9218 19071 9274 19080
rect 9126 19000 9182 19009
rect 9126 18935 9182 18944
rect 9140 18766 9168 18935
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9128 18624 9180 18630
rect 9126 18592 9128 18601
rect 9180 18592 9182 18601
rect 9126 18527 9182 18536
rect 9140 18426 9168 18527
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 9048 14521 9076 18362
rect 9232 17678 9260 19071
rect 9416 18698 9444 19858
rect 9508 19145 9536 22714
rect 9600 20534 9628 24142
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9692 23322 9720 24006
rect 10152 23798 10180 26200
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 22234 9812 23054
rect 9968 22710 9996 23258
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 10152 22030 10180 23190
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9876 21729 9904 21898
rect 9862 21720 9918 21729
rect 9862 21655 9918 21664
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 9954 20904 10010 20913
rect 9954 20839 10010 20848
rect 9968 20806 9996 20839
rect 10152 20806 10180 21286
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9494 19136 9550 19145
rect 9494 19071 9550 19080
rect 9586 19000 9642 19009
rect 9586 18935 9642 18944
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9600 18630 9628 18935
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9508 18465 9536 18566
rect 9494 18456 9550 18465
rect 9494 18391 9550 18400
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9416 17513 9444 18022
rect 9402 17504 9458 17513
rect 9402 17439 9458 17448
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9232 16250 9260 16662
rect 9310 16280 9366 16289
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9220 16244 9272 16250
rect 9310 16215 9366 16224
rect 9220 16186 9272 16192
rect 9140 15473 9168 16186
rect 9324 16114 9352 16215
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9126 15464 9182 15473
rect 9126 15399 9182 15408
rect 9034 14512 9090 14521
rect 9034 14447 9090 14456
rect 8758 14376 8814 14385
rect 8758 14311 8814 14320
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 9600 13326 9628 18226
rect 9692 17678 9720 18566
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9692 17270 9720 17614
rect 9784 17338 9812 19722
rect 10046 19680 10102 19689
rect 10046 19615 10102 19624
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9876 17338 9904 17478
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9968 16794 9996 18226
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9954 16688 10010 16697
rect 9954 16623 10010 16632
rect 9968 16454 9996 16623
rect 10060 16454 10088 19615
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10152 16046 10180 19994
rect 10244 16794 10272 24890
rect 10520 23186 10548 26200
rect 10888 23798 10916 26200
rect 10968 24268 11020 24274
rect 11072 24256 11100 26302
rect 11242 26200 11298 26302
rect 11610 26200 11666 27000
rect 11978 26330 12034 27000
rect 11978 26302 12296 26330
rect 11978 26200 12034 26302
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11020 24228 11100 24256
rect 10968 24210 11020 24216
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11152 22500 11204 22506
rect 11152 22442 11204 22448
rect 10508 22160 10560 22166
rect 10508 22102 10560 22108
rect 10520 21865 10548 22102
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10506 21856 10562 21865
rect 10506 21791 10562 21800
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10428 20874 10456 21354
rect 10612 20874 10640 21966
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10704 21010 10732 21286
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10600 20460 10652 20466
rect 10520 20420 10600 20448
rect 10322 19816 10378 19825
rect 10322 19751 10378 19760
rect 10336 19394 10364 19751
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 19514 10456 19654
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10336 19366 10456 19394
rect 10520 19378 10548 20420
rect 10600 20402 10652 20408
rect 10704 20398 10732 20946
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10600 19984 10652 19990
rect 10704 19961 10732 20198
rect 10796 20058 10824 20538
rect 10888 20466 10916 21558
rect 11164 21486 11192 22442
rect 11348 21962 11376 22646
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 21622 11376 21898
rect 11336 21616 11388 21622
rect 11336 21558 11388 21564
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10980 20942 11008 21286
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 11242 20904 11298 20913
rect 11242 20839 11298 20848
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10980 20074 11008 20402
rect 10784 20052 10836 20058
rect 10980 20046 11100 20074
rect 10784 19994 10836 20000
rect 10600 19926 10652 19932
rect 10690 19952 10746 19961
rect 10428 19242 10456 19366
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10520 18766 10548 19314
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10520 17338 10548 18702
rect 10612 18086 10640 19926
rect 10690 19887 10746 19896
rect 10876 19916 10928 19922
rect 10704 19310 10732 19887
rect 10876 19858 10928 19864
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10796 19174 10824 19654
rect 10888 19514 10916 19858
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10782 19000 10838 19009
rect 10782 18935 10838 18944
rect 10796 18222 10824 18935
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10428 17184 10456 17274
rect 10428 17156 10640 17184
rect 10612 17066 10640 17156
rect 10888 17134 10916 18566
rect 10980 17542 11008 19858
rect 11072 19786 11100 20046
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 11058 19408 11114 19417
rect 11058 19343 11114 19352
rect 11072 19242 11100 19343
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11058 18456 11114 18465
rect 11058 18391 11114 18400
rect 11072 18154 11100 18391
rect 11164 18358 11192 18770
rect 11256 18698 11284 20839
rect 11334 20768 11390 20777
rect 11334 20703 11390 20712
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17338 11008 17478
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11164 17270 11192 17614
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 11072 16794 11100 17138
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10244 16114 10272 16730
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10980 16250 11008 16594
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 16425 11100 16526
rect 11058 16416 11114 16425
rect 11058 16351 11114 16360
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11072 16182 11100 16351
rect 11348 16289 11376 20703
rect 11440 18290 11468 22578
rect 11532 21185 11560 24754
rect 11624 23186 11652 26200
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11900 23866 11928 24142
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 12268 23662 12296 26302
rect 12346 26200 12402 27000
rect 12714 26330 12770 27000
rect 12636 26302 12770 26330
rect 12360 24256 12388 26200
rect 12530 24304 12586 24313
rect 12440 24268 12492 24274
rect 12360 24228 12440 24256
rect 12530 24239 12586 24248
rect 12440 24210 12492 24216
rect 12544 24206 12572 24239
rect 12532 24200 12584 24206
rect 12438 24168 12494 24177
rect 12532 24142 12584 24148
rect 12438 24103 12494 24112
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11716 22982 11744 23054
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11978 22808 12034 22817
rect 11978 22743 12034 22752
rect 11888 22500 11940 22506
rect 11888 22442 11940 22448
rect 11900 22166 11928 22442
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11518 21176 11574 21185
rect 11518 21111 11574 21120
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11532 19446 11560 20470
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11900 19514 11928 19722
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11520 19440 11572 19446
rect 11520 19382 11572 19388
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11532 17814 11560 18634
rect 11624 18358 11652 18702
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11716 16674 11744 19314
rect 11992 18986 12020 22743
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 22098 12204 22510
rect 12268 22438 12296 22646
rect 12348 22568 12400 22574
rect 12348 22510 12400 22516
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12360 22273 12388 22510
rect 12346 22264 12402 22273
rect 12346 22199 12402 22208
rect 12254 22128 12310 22137
rect 12164 22092 12216 22098
rect 12452 22114 12480 24103
rect 12636 22710 12664 26302
rect 12714 26200 12770 26302
rect 13082 26200 13138 27000
rect 13450 26200 13506 27000
rect 13818 26200 13874 27000
rect 14186 26330 14242 27000
rect 14554 26330 14610 27000
rect 13924 26302 14242 26330
rect 13096 24596 13124 26200
rect 13464 24818 13492 26200
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 12820 24568 13124 24596
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12728 23497 12756 24278
rect 12714 23488 12770 23497
rect 12714 23423 12770 23432
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12624 22432 12676 22438
rect 12820 22409 12848 24568
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13740 23633 13768 24142
rect 13726 23624 13782 23633
rect 13726 23559 13782 23568
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13556 22642 13584 23122
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 12624 22374 12676 22380
rect 12806 22400 12862 22409
rect 12254 22063 12310 22072
rect 12360 22086 12480 22114
rect 12164 22034 12216 22040
rect 12070 21720 12126 21729
rect 12070 21655 12072 21664
rect 12124 21655 12126 21664
rect 12072 21626 12124 21632
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12176 20806 12204 21490
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12268 20602 12296 22063
rect 12360 20618 12388 22086
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21690 12480 21966
rect 12530 21720 12586 21729
rect 12440 21684 12492 21690
rect 12530 21655 12586 21664
rect 12440 21626 12492 21632
rect 12544 21570 12572 21655
rect 12452 21542 12572 21570
rect 12452 21350 12480 21542
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12544 21350 12572 21422
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12440 21072 12492 21078
rect 12438 21040 12440 21049
rect 12492 21040 12494 21049
rect 12438 20975 12494 20984
rect 12530 20768 12586 20777
rect 12452 20726 12530 20754
rect 12452 20618 12480 20726
rect 12530 20703 12586 20712
rect 12256 20596 12308 20602
rect 12360 20590 12480 20618
rect 12256 20538 12308 20544
rect 12636 20482 12664 22374
rect 12806 22335 12862 22344
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13268 22160 13320 22166
rect 13268 22102 13320 22108
rect 13280 21622 13308 22102
rect 13268 21616 13320 21622
rect 13268 21558 13320 21564
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12728 20942 12756 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 13372 20890 13400 22578
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 21593 13492 21830
rect 13450 21584 13506 21593
rect 13450 21519 13506 21528
rect 12452 20454 12664 20482
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11624 16646 11744 16674
rect 11808 18958 12020 18986
rect 11334 16280 11390 16289
rect 11334 16215 11390 16224
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10600 16040 10652 16046
rect 10968 16040 11020 16046
rect 10600 15982 10652 15988
rect 10966 16008 10968 16017
rect 11244 16040 11296 16046
rect 11020 16008 11022 16017
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10322 15600 10378 15609
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 10152 9042 10180 13126
rect 10244 10674 10272 15574
rect 10322 15535 10378 15544
rect 10336 15502 10364 15535
rect 10520 15502 10548 15982
rect 10612 15910 10640 15982
rect 11244 15982 11296 15988
rect 10966 15943 11022 15952
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10704 14958 10732 15438
rect 10966 15192 11022 15201
rect 11256 15162 11284 15982
rect 11532 15570 11560 16186
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 10966 15127 10968 15136
rect 11020 15127 11022 15136
rect 11244 15156 11296 15162
rect 10968 15098 11020 15104
rect 11244 15098 11296 15104
rect 10782 15056 10838 15065
rect 10782 14991 10784 15000
rect 10836 14991 10838 15000
rect 10784 14962 10836 14968
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14618 10640 14758
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10704 14414 10732 14894
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 13190 10732 14350
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 6840 2650 6868 8842
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 11624 6730 11652 16646
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16046 11744 16526
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11716 14958 11744 15982
rect 11808 15366 11836 18958
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11992 17746 12020 18770
rect 12084 18086 12112 19654
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12360 18834 12388 19314
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12268 18358 12296 18634
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12348 18216 12400 18222
rect 12176 18176 12348 18204
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11886 16280 11942 16289
rect 11886 16215 11942 16224
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11900 15094 11928 16215
rect 11992 15366 12020 17070
rect 12072 16448 12124 16454
rect 12176 16436 12204 18176
rect 12348 18158 12400 18164
rect 12348 17196 12400 17202
rect 12124 16408 12204 16436
rect 12268 17156 12348 17184
rect 12072 16390 12124 16396
rect 12084 16182 12112 16390
rect 12268 16182 12296 17156
rect 12348 17138 12400 17144
rect 12452 16538 12480 20454
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12530 19000 12586 19009
rect 12530 18935 12586 18944
rect 12544 18834 12572 18935
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 18154 12572 18226
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12636 17746 12664 20334
rect 12728 19378 12756 20878
rect 12820 20602 12848 20878
rect 13372 20862 13492 20890
rect 13360 20800 13412 20806
rect 12898 20768 12954 20777
rect 13360 20742 13412 20748
rect 12898 20703 12954 20712
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12912 20244 12940 20703
rect 12820 20216 12940 20244
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12728 17610 12756 18634
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 17202 12756 17546
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12452 16522 12572 16538
rect 12452 16516 12584 16522
rect 12452 16510 12532 16516
rect 12532 16458 12584 16464
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12440 16176 12492 16182
rect 12728 16164 12756 16458
rect 12492 16136 12756 16164
rect 12440 16118 12492 16124
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15638 12112 15982
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 12452 15450 12480 16118
rect 12360 15434 12480 15450
rect 12348 15428 12480 15434
rect 12400 15422 12480 15428
rect 12348 15370 12400 15376
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11992 14482 12020 15302
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 12084 13394 12112 15098
rect 12360 15042 12388 15370
rect 12440 15088 12492 15094
rect 12360 15036 12440 15042
rect 12360 15030 12492 15036
rect 12360 15014 12480 15030
rect 12360 14346 12388 15014
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14618 12480 14894
rect 12820 14618 12848 20216
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19990 13400 20742
rect 13464 20602 13492 20862
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13556 20466 13584 22578
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13648 21146 13676 22170
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13740 22030 13768 22102
rect 13832 22094 13860 26200
rect 13924 24750 13952 26302
rect 14186 26200 14242 26302
rect 14292 26302 14610 26330
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13924 23254 13952 24210
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22710 14136 22918
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13832 22066 13952 22094
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13464 19786 13492 20402
rect 13556 19922 13584 20402
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13648 19854 13676 20810
rect 13740 19990 13768 21286
rect 13832 20874 13860 21558
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13924 19854 13952 22066
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13268 19440 13320 19446
rect 13372 19428 13400 19722
rect 13452 19440 13504 19446
rect 13372 19400 13452 19428
rect 13268 19382 13320 19388
rect 13452 19382 13504 19388
rect 13280 19156 13308 19382
rect 13452 19168 13504 19174
rect 13280 19128 13400 19156
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 16998 13400 19128
rect 13450 19136 13452 19145
rect 13504 19136 13506 19145
rect 13450 19071 13506 19080
rect 13450 19000 13506 19009
rect 13450 18935 13506 18944
rect 13464 18834 13492 18935
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 17746 13492 18566
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13740 16658 13768 17750
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13818 17232 13874 17241
rect 13818 17167 13874 17176
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13832 15910 13860 17167
rect 13924 17134 13952 17546
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13174 15192 13230 15201
rect 13174 15127 13230 15136
rect 13188 14929 13216 15127
rect 13174 14920 13230 14929
rect 13174 14855 13230 14864
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14618 13400 15370
rect 13450 15056 13506 15065
rect 13450 14991 13506 15000
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12360 13138 12388 14282
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 14074 12756 14214
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12820 13938 12848 14554
rect 13464 14074 13492 14991
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 12440 13184 12492 13190
rect 12360 13132 12440 13138
rect 12360 13126 12492 13132
rect 12360 13110 12480 13126
rect 12360 8906 12388 13110
rect 13188 12918 13216 13466
rect 13740 13258 13768 15506
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13832 14006 13860 14554
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13924 13870 13952 15030
rect 14016 14550 14044 22102
rect 14096 21956 14148 21962
rect 14096 21898 14148 21904
rect 14108 21593 14136 21898
rect 14094 21584 14150 21593
rect 14094 21519 14150 21528
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14108 21010 14136 21286
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 14200 20210 14228 24754
rect 14292 24138 14320 26302
rect 14554 26200 14610 26302
rect 14922 26200 14978 27000
rect 15290 26330 15346 27000
rect 15212 26302 15346 26330
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14292 23730 14320 23802
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14292 22409 14320 22646
rect 14278 22400 14334 22409
rect 14278 22335 14334 22344
rect 14292 22012 14320 22335
rect 14384 22166 14412 24074
rect 14568 23905 14596 24074
rect 14554 23896 14610 23905
rect 14554 23831 14610 23840
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 14292 21984 14412 22012
rect 14278 21584 14334 21593
rect 14278 21519 14334 21528
rect 14292 21078 14320 21519
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14280 20868 14332 20874
rect 14384 20856 14412 21984
rect 14476 20942 14504 23054
rect 14568 22778 14596 23598
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14568 21690 14596 22714
rect 14752 22166 14780 24618
rect 14936 23322 14964 26200
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 15212 23202 15240 26302
rect 15290 26200 15346 26302
rect 15658 26330 15714 27000
rect 15658 26302 15884 26330
rect 15658 26200 15714 26302
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15488 24410 15516 24550
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15658 23352 15714 23361
rect 15658 23287 15714 23296
rect 14936 23174 15240 23202
rect 14740 22160 14792 22166
rect 14740 22102 14792 22108
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14332 20828 14412 20856
rect 14280 20810 14332 20816
rect 14292 20534 14320 20810
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14108 20182 14228 20210
rect 14108 19972 14136 20182
rect 14108 19944 14228 19972
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14108 16726 14136 18770
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14108 15026 14136 16050
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14200 14074 14228 19944
rect 14370 19952 14426 19961
rect 14280 19916 14332 19922
rect 14370 19887 14372 19896
rect 14280 19858 14332 19864
rect 14424 19887 14426 19896
rect 14372 19858 14424 19864
rect 14292 18766 14320 19858
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18426 14320 18702
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14292 17746 14320 18362
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14292 16658 14320 17682
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 14482 14320 15438
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14292 14006 14320 14418
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 14292 13394 14320 13942
rect 14384 13870 14412 19654
rect 14568 19514 14596 19790
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18630 14596 19110
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14660 16969 14688 21898
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 19009 14780 20742
rect 14936 20641 14964 23174
rect 15672 23050 15700 23287
rect 15476 23044 15528 23050
rect 15476 22986 15528 22992
rect 15660 23044 15712 23050
rect 15660 22986 15712 22992
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15120 22030 15148 22578
rect 15488 22098 15516 22986
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15028 21554 15056 21966
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15028 20942 15056 21286
rect 15212 21010 15240 22034
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 14922 20632 14978 20641
rect 14832 20596 14884 20602
rect 14922 20567 14978 20576
rect 14832 20538 14884 20544
rect 14844 19514 14872 20538
rect 15028 20398 15056 20878
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14830 19408 14886 19417
rect 14830 19343 14886 19352
rect 14738 19000 14794 19009
rect 14738 18935 14794 18944
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18222 14780 18566
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14646 16960 14702 16969
rect 14646 16895 14702 16904
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14568 16164 14596 16594
rect 14476 16136 14596 16164
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14476 13546 14504 16136
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 14346 14596 15982
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 14958 14688 15846
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14568 14074 14596 14282
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14384 13518 14504 13546
rect 14280 13388 14332 13394
rect 14200 13348 14280 13376
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12918 13676 13126
rect 14200 12986 14228 13348
rect 14280 13330 14332 13336
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14292 11626 14320 12174
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 14384 9178 14412 13518
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14660 12986 14688 13194
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14462 12608 14518 12617
rect 14462 12543 14518 12552
rect 14476 11898 14504 12543
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14568 11694 14596 12174
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 14752 8634 14780 17138
rect 14844 14278 14872 19343
rect 14936 18834 14964 20266
rect 15120 20262 15148 20946
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15212 20505 15240 20538
rect 15198 20496 15254 20505
rect 15198 20431 15254 20440
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15028 20058 15056 20198
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14922 18456 14978 18465
rect 14922 18391 14978 18400
rect 14936 16969 14964 18391
rect 15028 18290 15056 19382
rect 15120 19310 15148 20198
rect 15212 19689 15240 20334
rect 15304 19768 15332 21490
rect 15396 21418 15424 21898
rect 15474 21720 15530 21729
rect 15474 21655 15530 21664
rect 15488 21486 15516 21655
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15384 19780 15436 19786
rect 15304 19740 15384 19768
rect 15198 19680 15254 19689
rect 15198 19615 15254 19624
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15304 19174 15332 19740
rect 15384 19722 15436 19728
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15014 18048 15070 18057
rect 15014 17983 15070 17992
rect 14922 16960 14978 16969
rect 14922 16895 14978 16904
rect 15028 14618 15056 17983
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15120 15706 15148 17546
rect 15212 17082 15240 17546
rect 15304 17202 15332 19110
rect 15396 18970 15424 19246
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15488 18680 15516 20810
rect 15396 18652 15516 18680
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15212 17054 15332 17082
rect 15304 16522 15332 17054
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15304 15434 15332 16458
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 15304 14346 15332 15370
rect 15396 15162 15424 18652
rect 15580 18408 15608 22510
rect 15672 22409 15700 22986
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15658 22400 15714 22409
rect 15658 22335 15714 22344
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19446 15700 19858
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15488 18380 15608 18408
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15488 14958 15516 18380
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15580 18193 15608 18226
rect 15660 18216 15712 18222
rect 15566 18184 15622 18193
rect 15660 18158 15712 18164
rect 15566 18119 15622 18128
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15580 17610 15608 18022
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15672 16046 15700 18158
rect 15660 16040 15712 16046
rect 15566 16008 15622 16017
rect 15660 15982 15712 15988
rect 15566 15943 15568 15952
rect 15620 15943 15622 15952
rect 15568 15914 15620 15920
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15672 14618 15700 14962
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 15304 14006 15332 14282
rect 15764 14090 15792 22578
rect 15856 22506 15884 26302
rect 16026 26200 16082 27000
rect 16394 26330 16450 27000
rect 16224 26302 16450 26330
rect 16040 24682 16068 26200
rect 16118 24984 16174 24993
rect 16118 24919 16174 24928
rect 16028 24676 16080 24682
rect 16028 24618 16080 24624
rect 16132 24274 16160 24919
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 15948 23718 16160 23746
rect 15948 23186 15976 23718
rect 16132 23662 16160 23718
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 15934 22944 15990 22953
rect 15934 22879 15990 22888
rect 15948 22778 15976 22879
rect 15936 22772 15988 22778
rect 15936 22714 15988 22720
rect 15844 22500 15896 22506
rect 15844 22442 15896 22448
rect 16040 21690 16068 23598
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15856 18222 15884 18566
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15856 17202 15884 17818
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15856 16017 15884 16050
rect 15842 16008 15898 16017
rect 15842 15943 15898 15952
rect 15764 14074 15884 14090
rect 15764 14068 15896 14074
rect 15764 14062 15844 14068
rect 15844 14010 15896 14016
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15106 13424 15162 13433
rect 15106 13359 15162 13368
rect 15120 11898 15148 13359
rect 15304 13190 15332 13942
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15580 13462 15608 13670
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15842 12200 15898 12209
rect 15842 12135 15898 12144
rect 15856 11898 15884 12135
rect 15948 11898 15976 20402
rect 16040 19718 16068 21422
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18698 16068 19246
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 16040 16794 16068 18634
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16040 12170 16068 13738
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15856 11762 15884 11834
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 16132 9450 16160 21830
rect 16224 19378 16252 26302
rect 16394 26200 16450 26302
rect 16762 26200 16818 27000
rect 17130 26200 17186 27000
rect 17498 26330 17554 27000
rect 17498 26302 17632 26330
rect 17498 26200 17554 26302
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16408 24274 16436 24550
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16592 24070 16620 24686
rect 16776 24256 16804 26200
rect 17038 24848 17094 24857
rect 17038 24783 17094 24792
rect 16776 24228 16988 24256
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16316 23322 16344 23598
rect 16776 23497 16804 24074
rect 16762 23488 16818 23497
rect 16762 23423 16818 23432
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16762 22672 16818 22681
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16316 20398 16344 22510
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16408 22030 16436 22374
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16500 20992 16528 22646
rect 16762 22607 16818 22616
rect 16856 22636 16908 22642
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16592 21049 16620 22442
rect 16776 21894 16804 22607
rect 16856 22578 16908 22584
rect 16868 22506 16896 22578
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16960 22438 16988 24228
rect 17052 22778 17080 24783
rect 17144 23882 17172 26200
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17144 23854 17448 23882
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17144 22778 17172 23734
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 17328 23497 17356 23598
rect 17314 23488 17370 23497
rect 17314 23423 17370 23432
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17236 22642 17264 22918
rect 17420 22778 17448 23854
rect 17512 23662 17540 24074
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17604 23089 17632 26302
rect 17866 26200 17922 27000
rect 18234 26330 18290 27000
rect 18234 26302 18552 26330
rect 18234 26200 18290 26302
rect 17880 23882 17908 26200
rect 18524 24886 18552 26302
rect 18602 26200 18658 27000
rect 18970 26200 19026 27000
rect 19338 26200 19394 27000
rect 19706 26200 19762 27000
rect 20074 26330 20130 27000
rect 20166 26344 20222 26353
rect 20074 26302 20166 26330
rect 20074 26200 20130 26302
rect 20442 26330 20498 27000
rect 20166 26279 20222 26288
rect 20272 26302 20498 26330
rect 20272 26217 20300 26302
rect 20258 26208 20314 26217
rect 18512 24880 18564 24886
rect 18512 24822 18564 24828
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18524 24206 18552 24346
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17696 23854 17908 23882
rect 17590 23080 17646 23089
rect 17590 23015 17646 23024
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16854 21856 16910 21865
rect 16854 21791 16910 21800
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16408 20964 16528 20992
rect 16578 21040 16634 21049
rect 16578 20975 16634 20984
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16224 18086 16252 18634
rect 16316 18290 16344 19654
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16210 17912 16266 17921
rect 16210 17847 16266 17856
rect 16224 17649 16252 17847
rect 16210 17640 16266 17649
rect 16210 17575 16266 17584
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16224 16250 16252 17070
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 11762 16344 13126
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16408 11354 16436 20964
rect 16684 20806 16712 21286
rect 16868 21146 16896 21791
rect 17420 21690 17448 22034
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 16946 21312 17002 21321
rect 16946 21247 17002 21256
rect 16960 21146 16988 21247
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16762 20904 16818 20913
rect 16762 20839 16764 20848
rect 16816 20839 16818 20848
rect 16764 20810 16816 20816
rect 16672 20800 16724 20806
rect 16948 20800 17000 20806
rect 16672 20742 16724 20748
rect 16762 20768 16818 20777
rect 16948 20742 17000 20748
rect 16762 20703 16818 20712
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16500 19378 16528 20334
rect 16578 19952 16634 19961
rect 16578 19887 16634 19896
rect 16592 19446 16620 19887
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16500 18834 16528 19314
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16592 17882 16620 19246
rect 16670 19136 16726 19145
rect 16670 19071 16726 19080
rect 16684 18601 16712 19071
rect 16670 18592 16726 18601
rect 16670 18527 16726 18536
rect 16776 18057 16804 20703
rect 16854 20224 16910 20233
rect 16854 20159 16910 20168
rect 16762 18048 16818 18057
rect 16762 17983 16818 17992
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 17241 16528 17614
rect 16486 17232 16542 17241
rect 16486 17167 16542 17176
rect 16592 17082 16620 17682
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16500 17054 16620 17082
rect 16500 15570 16528 17054
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16500 14550 16528 15506
rect 16592 15366 16620 16934
rect 16684 16794 16712 17206
rect 16672 16788 16724 16794
rect 16868 16776 16896 20159
rect 16672 16730 16724 16736
rect 16776 16748 16896 16776
rect 16776 16289 16804 16748
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16762 16280 16818 16289
rect 16762 16215 16818 16224
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16776 15162 16804 15982
rect 16868 15162 16896 16594
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16868 15026 16896 15098
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16960 14906 16988 20742
rect 17052 19417 17080 21626
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17038 19408 17094 19417
rect 17038 19343 17094 19352
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17052 19009 17080 19110
rect 17038 19000 17094 19009
rect 17038 18935 17094 18944
rect 17144 18290 17172 20810
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17314 20360 17370 20369
rect 17236 18970 17264 20334
rect 17314 20295 17370 20304
rect 17328 19553 17356 20295
rect 17314 19544 17370 19553
rect 17314 19479 17370 19488
rect 17420 19417 17448 21490
rect 17512 21486 17540 22918
rect 17592 22500 17644 22506
rect 17696 22488 17724 23854
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 17868 23656 17920 23662
rect 18432 23633 18460 23734
rect 17868 23598 17920 23604
rect 18418 23624 18474 23633
rect 17880 23202 17908 23598
rect 18418 23559 18474 23568
rect 17958 23352 18014 23361
rect 17958 23287 18014 23296
rect 17644 22460 17724 22488
rect 17788 23186 17908 23202
rect 17788 23180 17920 23186
rect 17788 23174 17868 23180
rect 17592 22442 17644 22448
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 21690 17724 21830
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17788 21554 17816 23174
rect 17868 23122 17920 23128
rect 17972 23050 18000 23287
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18524 22778 18552 23190
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 18328 22500 18380 22506
rect 18328 22442 18380 22448
rect 17880 21962 17908 22442
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17696 20074 17724 21422
rect 17696 20058 17816 20074
rect 17696 20052 17828 20058
rect 17696 20046 17776 20052
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17406 19408 17462 19417
rect 17406 19343 17462 19352
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17052 17338 17080 17478
rect 17236 17338 17264 18090
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16726 17080 16934
rect 17040 16720 17092 16726
rect 17328 16697 17356 18362
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17420 17814 17448 18158
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17270 17448 17478
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17040 16662 17092 16668
rect 17314 16688 17370 16697
rect 17314 16623 17370 16632
rect 17316 16448 17368 16454
rect 17222 16416 17278 16425
rect 17316 16390 17368 16396
rect 17222 16351 17278 16360
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17038 16008 17094 16017
rect 17038 15943 17040 15952
rect 17092 15943 17094 15952
rect 17040 15914 17092 15920
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16776 14878 16988 14906
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16684 14346 16712 14826
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16500 13258 16528 13874
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12594 16528 13194
rect 16500 12566 16712 12594
rect 16684 12442 16712 12566
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 16592 11830 16620 12271
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16776 10810 16804 14878
rect 17052 14278 17080 15438
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16868 9110 16896 11562
rect 16960 11150 16988 13330
rect 17052 12646 17080 14214
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17052 12306 17080 12582
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11830 17080 12242
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 17144 4078 17172 16050
rect 17236 16017 17264 16351
rect 17222 16008 17278 16017
rect 17222 15943 17278 15952
rect 17328 15570 17356 16390
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17236 15094 17264 15302
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17328 14346 17356 15370
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17236 12434 17264 14010
rect 17328 13938 17356 14282
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17420 13530 17448 17070
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17236 12406 17448 12434
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17236 11830 17264 12310
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17328 10266 17356 10610
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17420 9654 17448 12406
rect 17512 10266 17540 19722
rect 17604 17338 17632 19722
rect 17696 19310 17724 20046
rect 17776 19994 17828 20000
rect 17880 19854 17908 21898
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18052 21412 18104 21418
rect 18052 21354 18104 21360
rect 18064 20806 18092 21354
rect 18340 20874 18368 22442
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17972 19854 18000 20198
rect 18326 20088 18382 20097
rect 18326 20023 18382 20032
rect 18340 19990 18368 20023
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17960 19712 18012 19718
rect 17880 19672 17960 19700
rect 17684 19304 17736 19310
rect 17880 19281 17908 19672
rect 17960 19654 18012 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 18050 19408 18106 19417
rect 17972 19310 18000 19382
rect 18050 19343 18106 19352
rect 17960 19304 18012 19310
rect 17684 19246 17736 19252
rect 17866 19272 17922 19281
rect 17960 19246 18012 19252
rect 17866 19207 17922 19216
rect 17972 18698 18000 19246
rect 18064 18766 18092 19343
rect 18432 18902 18460 22578
rect 18616 22234 18644 26200
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18696 23792 18748 23798
rect 18696 23734 18748 23740
rect 18708 23361 18736 23734
rect 18694 23352 18750 23361
rect 18694 23287 18750 23296
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18524 21486 18552 22034
rect 18694 21992 18750 22001
rect 18604 21956 18656 21962
rect 18694 21927 18750 21936
rect 18604 21898 18656 21904
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18524 20602 18552 21422
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18524 19310 18552 20402
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17604 14006 17632 16730
rect 17696 14074 17724 18566
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17788 15745 17816 17206
rect 17880 17202 17908 17478
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17880 16130 17908 16458
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17880 16114 18000 16130
rect 17880 16108 18012 16114
rect 17880 16102 17960 16108
rect 17960 16050 18012 16056
rect 17774 15736 17830 15745
rect 17774 15671 17830 15680
rect 17776 15428 17828 15434
rect 17972 15416 18000 16050
rect 17828 15388 18000 15416
rect 17776 15370 17828 15376
rect 17788 15094 17816 15370
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 18340 14550 18368 18770
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18432 17202 18460 18362
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18524 16250 18552 18294
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18524 14346 18552 16186
rect 18616 14906 18644 21898
rect 18708 21894 18736 21927
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18800 21706 18828 24822
rect 18984 24721 19012 26200
rect 18970 24712 19026 24721
rect 18970 24647 19026 24656
rect 19352 24313 19380 26200
rect 19338 24304 19394 24313
rect 19156 24268 19208 24274
rect 19338 24239 19394 24248
rect 19156 24210 19208 24216
rect 19168 23662 19196 24210
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19246 23624 19302 23633
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 18892 22778 18920 23462
rect 19168 23322 19196 23598
rect 19246 23559 19248 23568
rect 19300 23559 19302 23568
rect 19248 23530 19300 23536
rect 19246 23352 19302 23361
rect 19156 23316 19208 23322
rect 19246 23287 19302 23296
rect 19156 23258 19208 23264
rect 19260 23050 19288 23287
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 19156 22704 19208 22710
rect 19156 22646 19208 22652
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18892 21865 18920 22170
rect 18878 21856 18934 21865
rect 18878 21791 18934 21800
rect 18800 21678 19104 21706
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18800 21010 18828 21558
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 21078 18920 21422
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 17882 18736 20742
rect 18800 20466 18828 20946
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18970 19272 19026 19281
rect 18970 19207 19026 19216
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16114 18736 16458
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18800 15706 18828 18906
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18800 14958 18828 15642
rect 18788 14952 18840 14958
rect 18616 14878 18736 14906
rect 18788 14894 18840 14900
rect 18892 14890 18920 18838
rect 18984 16250 19012 19207
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14482 18644 14758
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 18524 14006 18552 14282
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 17592 13864 17644 13870
rect 17776 13864 17828 13870
rect 17644 13812 17776 13818
rect 17592 13806 17828 13812
rect 17604 13790 17816 13806
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12918 18368 13942
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17880 11801 17908 12786
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18248 12322 18276 12718
rect 18432 12442 18460 13874
rect 18708 13818 18736 14878
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18524 13790 18736 13818
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18248 12294 18460 12322
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18144 11824 18196 11830
rect 17866 11792 17922 11801
rect 18340 11778 18368 12174
rect 18196 11772 18368 11778
rect 18144 11766 18368 11772
rect 17866 11727 17922 11736
rect 18156 11750 18368 11766
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17590 11248 17646 11257
rect 17590 11183 17646 11192
rect 17604 10742 17632 11183
rect 17696 11082 17724 11494
rect 18156 11082 18184 11750
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18432 11014 18460 12294
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18524 10810 18552 13790
rect 18694 13560 18750 13569
rect 18694 13495 18750 13504
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 17592 10736 17644 10742
rect 17960 10736 18012 10742
rect 17592 10678 17644 10684
rect 17788 10684 17960 10690
rect 17788 10678 18012 10684
rect 17788 10674 18000 10678
rect 18616 10674 18644 12582
rect 17776 10668 18000 10674
rect 17828 10662 18000 10668
rect 18604 10668 18656 10674
rect 17776 10610 17828 10616
rect 18604 10610 18656 10616
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 18050 9616 18106 9625
rect 18708 9586 18736 13495
rect 18800 12918 18828 14486
rect 18878 13696 18934 13705
rect 18878 13631 18934 13640
rect 18892 13530 18920 13631
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18984 13258 19012 15846
rect 19076 14278 19104 21678
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 19076 11812 19104 13942
rect 19168 13394 19196 22646
rect 19260 22080 19288 22986
rect 19352 22817 19380 24006
rect 19338 22808 19394 22817
rect 19338 22743 19394 22752
rect 19444 22681 19472 24006
rect 19720 23594 19748 26200
rect 20442 26200 20498 26302
rect 20810 26200 20866 27000
rect 21178 26330 21234 27000
rect 20916 26302 21234 26330
rect 20258 26143 20314 26152
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20732 24342 20760 24890
rect 19800 24336 19852 24342
rect 19800 24278 19852 24284
rect 20720 24336 20772 24342
rect 20720 24278 20772 24284
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19812 23526 19840 24278
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19628 23100 19656 23462
rect 19536 23072 19656 23100
rect 19904 23089 19932 24006
rect 20168 23588 20220 23594
rect 20168 23530 20220 23536
rect 19890 23080 19946 23089
rect 19536 22982 19564 23072
rect 19708 23044 19760 23050
rect 19890 23015 19946 23024
rect 19984 23044 20036 23050
rect 19708 22986 19760 22992
rect 19984 22986 20036 22992
rect 19524 22976 19576 22982
rect 19616 22976 19668 22982
rect 19524 22918 19576 22924
rect 19614 22944 19616 22953
rect 19668 22944 19670 22953
rect 19430 22672 19486 22681
rect 19430 22607 19486 22616
rect 19536 22574 19564 22918
rect 19727 22930 19755 22986
rect 19996 22953 20024 22986
rect 19982 22944 20038 22953
rect 19727 22902 19840 22930
rect 19614 22879 19670 22888
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19260 22052 19380 22080
rect 19352 20874 19380 22052
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19260 18834 19288 20402
rect 19444 20097 19472 22510
rect 19812 22506 19840 22902
rect 19982 22879 20038 22888
rect 19982 22808 20038 22817
rect 19982 22743 19984 22752
rect 20036 22743 20038 22752
rect 19984 22714 20036 22720
rect 19800 22500 19852 22506
rect 19800 22442 19852 22448
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 20777 19564 22374
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19628 20874 19656 21490
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19522 20768 19578 20777
rect 19522 20703 19578 20712
rect 19628 20534 19656 20810
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19430 20088 19486 20097
rect 19430 20023 19486 20032
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19514 19472 19654
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19432 19372 19484 19378
rect 19536 19360 19564 20334
rect 19720 19786 19748 21830
rect 19996 21690 20024 22442
rect 20076 22432 20128 22438
rect 20074 22400 20076 22409
rect 20128 22400 20130 22409
rect 20074 22335 20130 22344
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19890 21040 19946 21049
rect 19890 20975 19946 20984
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19812 19854 19840 20878
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 19484 19332 19564 19360
rect 19616 19372 19668 19378
rect 19432 19314 19484 19320
rect 19616 19314 19668 19320
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19352 18873 19380 19178
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19338 18864 19394 18873
rect 19248 18828 19300 18834
rect 19338 18799 19394 18808
rect 19248 18770 19300 18776
rect 19260 18426 19288 18770
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 16425 19288 17614
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19352 16658 19380 17274
rect 19430 16824 19486 16833
rect 19430 16759 19432 16768
rect 19484 16759 19486 16768
rect 19432 16730 19484 16736
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19246 16416 19302 16425
rect 19246 16351 19302 16360
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 18800 11784 19104 11812
rect 18050 9551 18106 9560
rect 18696 9580 18748 9586
rect 18064 9382 18092 9551
rect 18696 9522 18748 9528
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 9042 18736 9318
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18800 3058 18828 11784
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10810 18920 10950
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 19168 9674 19196 13194
rect 19260 11898 19288 16186
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19444 14074 19472 14962
rect 19536 14278 19564 19110
rect 19628 17921 19656 19314
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18970 19748 19246
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19904 18766 19932 20975
rect 20088 20262 20116 22034
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19614 17912 19670 17921
rect 19614 17847 19670 17856
rect 19798 17912 19854 17921
rect 19798 17847 19854 17856
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19444 13394 19472 14010
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19444 12986 19472 13330
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19444 12238 19472 12922
rect 19524 12436 19576 12442
rect 19628 12434 19656 17682
rect 19812 17542 19840 17847
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19720 15042 19748 17478
rect 19798 16688 19854 16697
rect 19798 16623 19854 16632
rect 19812 15434 19840 16623
rect 19904 16250 19932 18226
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19996 15722 20024 19654
rect 20180 19145 20208 23530
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20258 22808 20314 22817
rect 20258 22743 20314 22752
rect 20272 22710 20300 22743
rect 20260 22704 20312 22710
rect 20260 22646 20312 22652
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20272 21078 20300 21626
rect 20260 21072 20312 21078
rect 20260 21014 20312 21020
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 20058 20300 20198
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20166 19136 20222 19145
rect 20166 19071 20222 19080
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 17338 20208 18566
rect 20364 18222 20392 23462
rect 20456 22710 20484 24142
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20352 17264 20404 17270
rect 20350 17232 20352 17241
rect 20404 17232 20406 17241
rect 20168 17196 20220 17202
rect 20350 17167 20406 17176
rect 20168 17138 20220 17144
rect 20180 16522 20208 17138
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20456 16182 20484 21286
rect 20548 20641 20576 22578
rect 20626 22264 20682 22273
rect 20824 22234 20852 26200
rect 20626 22199 20682 22208
rect 20812 22228 20864 22234
rect 20640 20806 20668 22199
rect 20812 22170 20864 22176
rect 20718 21584 20774 21593
rect 20718 21519 20774 21528
rect 20812 21548 20864 21554
rect 20732 21010 20760 21519
rect 20812 21490 20864 21496
rect 20824 21457 20852 21490
rect 20810 21448 20866 21457
rect 20810 21383 20866 21392
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20534 20632 20590 20641
rect 20534 20567 20590 20576
rect 20732 20398 20760 20946
rect 20824 20602 20852 21082
rect 20916 20913 20944 26302
rect 21178 26200 21234 26302
rect 21456 26308 21508 26314
rect 21456 26250 21508 26256
rect 21468 26058 21496 26250
rect 21546 26200 21602 27000
rect 21914 26330 21970 27000
rect 21652 26302 21970 26330
rect 22192 26376 22244 26382
rect 22282 26330 22338 27000
rect 22650 26330 22706 27000
rect 23018 26330 23074 27000
rect 23386 26330 23442 27000
rect 22244 26324 22338 26330
rect 22192 26318 22338 26324
rect 22204 26302 22338 26318
rect 21560 26058 21588 26200
rect 21468 26030 21588 26058
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 21100 24206 21128 24686
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 21178 23216 21234 23225
rect 21178 23151 21234 23160
rect 20996 22432 21048 22438
rect 21192 22409 21220 23151
rect 20996 22374 21048 22380
rect 21178 22400 21234 22409
rect 21008 22137 21036 22374
rect 21178 22335 21234 22344
rect 20994 22128 21050 22137
rect 20994 22063 21050 22072
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21008 21350 21036 21898
rect 21284 21570 21312 23598
rect 21376 21894 21404 24142
rect 21456 23248 21508 23254
rect 21456 23190 21508 23196
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21192 21542 21312 21570
rect 21376 21554 21404 21830
rect 21364 21548 21416 21554
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 20902 20904 20958 20913
rect 20902 20839 20958 20848
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 20994 20768 21050 20777
rect 20994 20703 21050 20712
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20548 19446 20576 20266
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20626 19408 20682 19417
rect 20444 16176 20496 16182
rect 20444 16118 20496 16124
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19904 15694 20024 15722
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19904 15366 19932 15694
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19720 15014 19840 15042
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 13802 19748 14894
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19812 12986 19840 15014
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19904 12866 19932 14350
rect 19812 12838 19932 12866
rect 19576 12406 19656 12434
rect 19708 12436 19760 12442
rect 19524 12378 19576 12384
rect 19708 12378 19760 12384
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19260 10674 19288 11834
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 18984 9646 19196 9674
rect 18984 9586 19012 9646
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 19352 3058 19380 12106
rect 19444 11218 19472 12174
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19628 11830 19656 12038
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19720 11286 19748 12378
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19812 10674 19840 12838
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19996 10538 20024 15574
rect 20088 13530 20116 15982
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20088 12152 20116 12854
rect 20180 12714 20208 13670
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 20168 12164 20220 12170
rect 20088 12124 20168 12152
rect 20088 11830 20116 12124
rect 20168 12106 20220 12112
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 20272 11694 20300 15506
rect 20548 15502 20576 19382
rect 20626 19343 20628 19352
rect 20680 19343 20682 19352
rect 20628 19314 20680 19320
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 13394 20392 13670
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20088 11218 20116 11630
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20074 11112 20130 11121
rect 20074 11047 20130 11056
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19444 7886 19472 10406
rect 19522 10296 19578 10305
rect 20088 10266 20116 11047
rect 20180 10606 20208 11154
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19522 10231 19524 10240
rect 19576 10231 19578 10240
rect 20076 10260 20128 10266
rect 19524 10202 19576 10208
rect 20076 10202 20128 10208
rect 20088 10062 20116 10202
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19536 9178 19564 9522
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6748 800 6776 2382
rect 19536 2378 19564 2926
rect 20088 2446 20116 9658
rect 20180 9586 20208 10406
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20272 9382 20300 10066
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20364 8566 20392 12582
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20456 8498 20484 12582
rect 20548 10674 20576 13330
rect 20640 12288 20668 18022
rect 20732 13938 20760 19450
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20824 18737 20852 19246
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20810 18728 20866 18737
rect 20810 18663 20866 18672
rect 20916 18426 20944 19110
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20902 18320 20958 18329
rect 20902 18255 20904 18264
rect 20956 18255 20958 18264
rect 20904 18226 20956 18232
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20824 17338 20852 17546
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20810 17232 20866 17241
rect 20916 17218 20944 17546
rect 21008 17270 21036 20703
rect 21100 20534 21128 20810
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21100 19718 21128 20470
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 18698 21128 19654
rect 21192 19174 21220 21542
rect 21364 21490 21416 21496
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21178 19000 21234 19009
rect 21178 18935 21234 18944
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21192 18329 21220 18935
rect 21178 18320 21234 18329
rect 21178 18255 21234 18264
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20866 17190 20944 17218
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20810 17167 20866 17176
rect 20824 16572 20852 17167
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21008 16794 21036 17070
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20824 16544 20944 16572
rect 20810 15736 20866 15745
rect 20810 15671 20866 15680
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20824 12866 20852 15671
rect 20916 15076 20944 16544
rect 21008 16114 21036 16730
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20996 15088 21048 15094
rect 20916 15048 20996 15076
rect 20996 15030 21048 15036
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 14006 20944 14282
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20732 12838 20852 12866
rect 20732 12481 20760 12838
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20718 12472 20774 12481
rect 20718 12407 20774 12416
rect 20720 12300 20772 12306
rect 20640 12260 20720 12288
rect 20720 12242 20772 12248
rect 20824 12186 20852 12650
rect 21008 12628 21036 14010
rect 20732 12158 20852 12186
rect 20916 12600 21036 12628
rect 20732 11914 20760 12158
rect 20640 11886 20760 11914
rect 20640 11558 20668 11886
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20718 11520 20774 11529
rect 20718 11455 20774 11464
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20548 9722 20576 9998
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19524 2372 19576 2378
rect 19524 2314 19576 2320
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 800 20208 4014
rect 20640 3534 20668 11018
rect 20732 10198 20760 11455
rect 20810 11112 20866 11121
rect 20810 11047 20866 11056
rect 20824 10742 20852 11047
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 20916 10674 20944 12600
rect 20994 12472 21050 12481
rect 21100 12442 21128 18158
rect 21284 17728 21312 21422
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21376 17882 21404 19722
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21284 17700 21404 17728
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 15434 21220 16934
rect 21376 16726 21404 17700
rect 21468 17202 21496 23190
rect 21652 23066 21680 26302
rect 21914 26200 21970 26302
rect 22282 26200 22338 26302
rect 22388 26302 22706 26330
rect 21914 25664 21970 25673
rect 21914 25599 21970 25608
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21836 23186 21864 24346
rect 21928 24274 21956 25599
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 22020 23730 22048 24618
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22008 23316 22060 23322
rect 22112 23304 22140 23598
rect 22060 23276 22140 23304
rect 22008 23258 22060 23264
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21560 23038 21680 23066
rect 21916 23044 21968 23050
rect 21560 21185 21588 23038
rect 21916 22986 21968 22992
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21546 21176 21602 21185
rect 21546 21111 21602 21120
rect 21546 18728 21602 18737
rect 21546 18663 21602 18672
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21560 17105 21588 18663
rect 21546 17096 21602 17105
rect 21546 17031 21602 17040
rect 21364 16720 21416 16726
rect 21364 16662 21416 16668
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15570 21312 16390
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21376 15162 21404 16662
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 20994 12407 21050 12416
rect 21088 12436 21140 12442
rect 21008 11354 21036 12407
rect 21192 12434 21220 14486
rect 21284 13258 21312 15030
rect 21468 13954 21496 16390
rect 21652 16114 21680 22918
rect 21744 22438 21772 22918
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21744 21962 21772 22170
rect 21732 21956 21784 21962
rect 21732 21898 21784 21904
rect 21744 21078 21772 21898
rect 21732 21072 21784 21078
rect 21732 21014 21784 21020
rect 21836 19378 21864 22578
rect 21928 22234 21956 22986
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22020 22778 22048 22918
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 22020 22273 22048 22374
rect 22006 22264 22062 22273
rect 21916 22228 21968 22234
rect 22006 22199 22062 22208
rect 21916 22170 21968 22176
rect 21914 22128 21970 22137
rect 22112 22098 22140 23276
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 22296 23186 22324 23258
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22284 22772 22336 22778
rect 22388 22760 22416 26302
rect 22650 26200 22706 26302
rect 22756 26302 23074 26330
rect 22466 26072 22522 26081
rect 22466 26007 22522 26016
rect 22480 23798 22508 26007
rect 22560 24132 22612 24138
rect 22560 24074 22612 24080
rect 22468 23792 22520 23798
rect 22468 23734 22520 23740
rect 22468 23656 22520 23662
rect 22572 23610 22600 24074
rect 22520 23604 22600 23610
rect 22468 23598 22600 23604
rect 22336 22732 22416 22760
rect 22480 23582 22600 23598
rect 22284 22714 22336 22720
rect 22480 22658 22508 23582
rect 22756 22760 22784 26302
rect 23018 26200 23074 26302
rect 23308 26302 23442 26330
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22848 23798 22876 24074
rect 22836 23792 22888 23798
rect 22836 23734 22888 23740
rect 22848 22982 22876 23734
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23204 23248 23256 23254
rect 23204 23190 23256 23196
rect 23112 23044 23164 23050
rect 23112 22986 23164 22992
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22388 22630 22508 22658
rect 22572 22732 22784 22760
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 21914 22063 21970 22072
rect 22100 22092 22152 22098
rect 21928 21457 21956 22063
rect 22100 22034 22152 22040
rect 22112 21486 22140 22034
rect 22100 21480 22152 21486
rect 21914 21448 21970 21457
rect 22100 21422 22152 21428
rect 21914 21383 21970 21392
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22020 21078 22048 21286
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21928 19281 21956 20946
rect 22112 20942 22140 21422
rect 22204 21010 22232 22374
rect 22296 22166 22324 22442
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22388 22098 22416 22630
rect 22468 22568 22520 22574
rect 22468 22510 22520 22516
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22282 21992 22338 22001
rect 22282 21927 22338 21936
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22190 20904 22246 20913
rect 22112 19922 22140 20878
rect 22190 20839 22246 20848
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22008 19304 22060 19310
rect 21914 19272 21970 19281
rect 22008 19246 22060 19252
rect 21914 19207 21970 19216
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21928 17066 21956 17818
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21376 13926 21496 13954
rect 21376 13734 21404 13926
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13258 21404 13670
rect 21468 13530 21496 13738
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21284 12918 21312 13194
rect 21560 13190 21588 13738
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21272 12912 21324 12918
rect 21270 12880 21272 12889
rect 21324 12880 21326 12889
rect 21270 12815 21326 12824
rect 21364 12436 21416 12442
rect 21192 12406 21312 12434
rect 21088 12378 21140 12384
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21100 12102 21128 12242
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 21192 11898 21220 12174
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21086 11792 21142 11801
rect 21086 11727 21142 11736
rect 21100 11558 21128 11727
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 21192 10130 21220 11834
rect 21284 11150 21312 12406
rect 21364 12378 21416 12384
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21376 10554 21404 12378
rect 21652 12186 21680 15846
rect 21744 15366 21772 16934
rect 21836 16697 21864 16934
rect 21822 16688 21878 16697
rect 21822 16623 21878 16632
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21836 16250 21864 16526
rect 22020 16454 22048 19246
rect 22112 18086 22140 19858
rect 22204 18714 22232 20839
rect 22296 19145 22324 21927
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 21146 22416 21286
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22480 20505 22508 22510
rect 22572 22506 22600 22732
rect 22742 22672 22798 22681
rect 22742 22607 22798 22616
rect 22560 22500 22612 22506
rect 22560 22442 22612 22448
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 22664 21486 22692 21558
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22466 20496 22522 20505
rect 22466 20431 22522 20440
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22388 19514 22416 20198
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22480 19258 22508 20334
rect 22572 19514 22600 21422
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22664 19922 22692 20810
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22650 19816 22706 19825
rect 22650 19751 22706 19760
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22480 19230 22600 19258
rect 22468 19168 22520 19174
rect 22282 19136 22338 19145
rect 22468 19110 22520 19116
rect 22282 19071 22338 19080
rect 22204 18686 22416 18714
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22112 17746 22140 18022
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 22112 17202 22140 17682
rect 22192 17536 22244 17542
rect 22190 17504 22192 17513
rect 22244 17504 22246 17513
rect 22190 17439 22246 17448
rect 22296 17338 22324 18566
rect 22388 17338 22416 18686
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22006 16280 22062 16289
rect 21824 16244 21876 16250
rect 22006 16215 22008 16224
rect 21824 16186 21876 16192
rect 22060 16215 22062 16224
rect 22008 16186 22060 16192
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21916 14952 21968 14958
rect 22112 14940 22140 16594
rect 22296 16046 22324 17274
rect 22480 16969 22508 19110
rect 22572 18766 22600 19230
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22466 16960 22522 16969
rect 22466 16895 22522 16904
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 21968 14912 22140 14940
rect 21916 14894 21968 14900
rect 21928 14278 21956 14894
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21822 13968 21878 13977
rect 21822 13903 21878 13912
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21744 12442 21772 13670
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21652 12158 21772 12186
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21284 10526 21404 10554
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 9722 20760 9930
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 8566 20760 8774
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20824 5302 20852 8910
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 21284 4162 21312 10526
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21376 6798 21404 10406
rect 21468 7410 21496 12038
rect 21652 11762 21680 12038
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21548 11688 21600 11694
rect 21744 11642 21772 12158
rect 21548 11630 21600 11636
rect 21560 10130 21588 11630
rect 21652 11614 21772 11642
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21546 9616 21602 9625
rect 21546 9551 21602 9560
rect 21560 7886 21588 9551
rect 21652 7954 21680 11614
rect 21836 11150 21864 13903
rect 21928 13870 21956 14214
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21928 13326 21956 13806
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 13433 22232 13738
rect 22190 13424 22246 13433
rect 22190 13359 22246 13368
rect 21916 13320 21968 13326
rect 21968 13268 22048 13274
rect 21916 13262 22048 13268
rect 21928 13246 22048 13262
rect 22020 12782 22048 13246
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22204 12986 22232 13194
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 22020 12238 22048 12718
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21744 8498 21772 11018
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21836 9722 21864 9930
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21928 8022 21956 11630
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22020 11014 22048 11290
rect 22296 11098 22324 15438
rect 22112 11070 22324 11098
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 22112 5234 22140 11070
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22204 5710 22232 10066
rect 22296 6798 22324 10406
rect 22388 9518 22416 15846
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22480 15450 22508 15642
rect 22572 15638 22600 18566
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22480 15422 22600 15450
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22480 8106 22508 14826
rect 22572 8974 22600 15422
rect 22664 15094 22692 19751
rect 22756 18714 22784 22607
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 19990 22876 22510
rect 23124 22438 23152 22986
rect 23112 22432 23164 22438
rect 23216 22420 23244 23190
rect 23308 22545 23336 26302
rect 23386 26200 23442 26302
rect 24490 26200 24546 27000
rect 24858 26200 24914 27000
rect 24950 26480 25006 26489
rect 24950 26415 25006 26424
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23400 24041 23428 24754
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23386 24032 23442 24041
rect 23386 23967 23442 23976
rect 23860 23662 23888 24074
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23294 22536 23350 22545
rect 23294 22471 23350 22480
rect 23216 22392 23336 22420
rect 23112 22374 23164 22380
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22166 23336 22392
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 20602 23336 21966
rect 23400 21162 23428 22918
rect 23664 22432 23716 22438
rect 23662 22400 23664 22409
rect 23860 22420 23888 23598
rect 23716 22400 23718 22409
rect 23662 22335 23718 22344
rect 23768 22392 23888 22420
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23492 21894 23520 22102
rect 23768 22094 23796 22392
rect 23676 22066 23796 22094
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23584 21690 23612 21830
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23676 21350 23704 22066
rect 23848 21616 23900 21622
rect 23848 21558 23900 21564
rect 23756 21412 23808 21418
rect 23756 21354 23808 21360
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23400 21134 23612 21162
rect 23768 21146 23796 21354
rect 23400 21010 23428 21134
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23388 20800 23440 20806
rect 23386 20768 23388 20777
rect 23440 20768 23442 20777
rect 23386 20703 23442 20712
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23204 20528 23256 20534
rect 23202 20496 23204 20505
rect 23256 20496 23258 20505
rect 23202 20431 23258 20440
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22848 18834 22876 19926
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22756 18686 22876 18714
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22756 18057 22784 18362
rect 22848 18222 22876 18686
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22940 18358 22968 18566
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22742 18048 22798 18057
rect 22742 17983 22798 17992
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17785 23336 19654
rect 23400 19310 23428 20334
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23400 18086 23428 19246
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23386 17912 23442 17921
rect 23386 17847 23388 17856
rect 23440 17847 23442 17856
rect 23388 17818 23440 17824
rect 23294 17776 23350 17785
rect 23492 17746 23520 20946
rect 23584 18086 23612 21134
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23860 20942 23888 21558
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23294 17711 23350 17720
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23386 17640 23442 17649
rect 23386 17575 23388 17584
rect 23440 17575 23442 17584
rect 23388 17546 23440 17552
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22756 14940 22784 17478
rect 23492 17354 23520 17682
rect 23296 17332 23348 17338
rect 23492 17326 23612 17354
rect 23296 17274 23348 17280
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 15892 23336 17274
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23386 17096 23442 17105
rect 23386 17031 23442 17040
rect 23400 16017 23428 17031
rect 23492 16504 23520 17138
rect 23584 16658 23612 17326
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23572 16516 23624 16522
rect 23492 16476 23572 16504
rect 23572 16458 23624 16464
rect 23386 16008 23442 16017
rect 23386 15943 23442 15952
rect 23308 15864 23428 15892
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 22664 14912 22784 14940
rect 22664 13705 22692 14912
rect 22742 13968 22798 13977
rect 22742 13903 22798 13912
rect 22650 13696 22706 13705
rect 22650 13631 22706 13640
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22664 12889 22692 13194
rect 22650 12880 22706 12889
rect 22650 12815 22706 12824
rect 22664 12170 22692 12815
rect 22652 12164 22704 12170
rect 22652 12106 22704 12112
rect 22664 10062 22692 12106
rect 22756 10470 22784 13903
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22388 8078 22508 8106
rect 22664 8090 22692 8910
rect 22652 8084 22704 8090
rect 22388 6914 22416 8078
rect 22652 8026 22704 8032
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22388 6886 22508 6914
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22480 4622 22508 6886
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 21192 4146 21312 4162
rect 21180 4140 21312 4146
rect 21232 4134 21312 4140
rect 21180 4082 21232 4088
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22020 1170 22048 3402
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 22112 2009 22140 2314
rect 22098 2000 22154 2009
rect 22098 1935 22154 1944
rect 22204 1601 22232 4014
rect 22756 3602 22784 7142
rect 22848 4146 22876 15302
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23018 13016 23074 13025
rect 23018 12951 23074 12960
rect 22928 12912 22980 12918
rect 22926 12880 22928 12889
rect 22980 12880 22982 12889
rect 22926 12815 22982 12824
rect 23032 12646 23060 12951
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11082 23336 15302
rect 23400 14770 23428 15864
rect 23584 15076 23612 16458
rect 23676 15502 23704 19382
rect 23846 18864 23902 18873
rect 23846 18799 23848 18808
rect 23900 18799 23902 18808
rect 23848 18770 23900 18776
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23860 17338 23888 17682
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23952 17066 23980 24006
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 24044 23050 24072 23258
rect 24032 23044 24084 23050
rect 24032 22986 24084 22992
rect 24044 21690 24072 22986
rect 24122 21992 24178 22001
rect 24122 21927 24178 21936
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24136 21049 24164 21927
rect 24228 21146 24256 24550
rect 24504 24206 24532 26200
rect 24766 25256 24822 25265
rect 24766 25191 24822 25200
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24780 23798 24808 25191
rect 24768 23792 24820 23798
rect 24768 23734 24820 23740
rect 24964 23254 24992 26415
rect 25226 26200 25282 27000
rect 25044 24064 25096 24070
rect 25044 24006 25096 24012
rect 25056 23866 25084 24006
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 24952 23248 25004 23254
rect 24952 23190 25004 23196
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24504 22166 24532 22578
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24492 22160 24544 22166
rect 24492 22102 24544 22108
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24122 21040 24178 21049
rect 24122 20975 24178 20984
rect 24030 20904 24086 20913
rect 24030 20839 24032 20848
rect 24084 20839 24086 20848
rect 24032 20810 24084 20816
rect 24228 20398 24256 21082
rect 24504 20942 24532 22102
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24320 20534 24348 20878
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24308 20528 24360 20534
rect 24308 20470 24360 20476
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24320 19854 24348 20470
rect 24308 19848 24360 19854
rect 24308 19790 24360 19796
rect 24320 19446 24348 19790
rect 24308 19440 24360 19446
rect 24308 19382 24360 19388
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 23940 17060 23992 17066
rect 23940 17002 23992 17008
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23664 15088 23716 15094
rect 23584 15048 23664 15076
rect 23664 15030 23716 15036
rect 23400 14742 23520 14770
rect 23386 14648 23442 14657
rect 23386 14583 23388 14592
rect 23440 14583 23442 14592
rect 23388 14554 23440 14560
rect 23492 14498 23520 14742
rect 23400 14470 23520 14498
rect 23400 11665 23428 14470
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23584 14074 23612 14282
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23492 12782 23520 14010
rect 23676 13938 23704 15030
rect 23768 14521 23796 16934
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23952 16046 23980 16390
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23952 14958 23980 15982
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 24044 14634 24072 18770
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 23952 14606 24072 14634
rect 23754 14512 23810 14521
rect 23754 14447 23810 14456
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23386 11656 23442 11665
rect 23386 11591 23442 11600
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 23032 9722 23060 9862
rect 23294 9752 23350 9761
rect 23020 9716 23072 9722
rect 23294 9687 23350 9696
rect 23020 9658 23072 9664
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 7410 23428 9318
rect 23492 8634 23520 11698
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23584 8022 23612 13194
rect 23676 12889 23704 13874
rect 23662 12880 23718 12889
rect 23662 12815 23718 12824
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22296 3058 22324 3334
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 2446 23336 5782
rect 23860 3058 23888 14214
rect 23952 12714 23980 14606
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24044 13870 24072 14418
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 24044 12306 24072 13806
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23952 10674 23980 11290
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23952 9586 23980 9930
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24044 8922 24072 11222
rect 24136 10062 24164 18566
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24228 12442 24256 16050
rect 24320 15178 24348 17478
rect 24412 16250 24440 20742
rect 24492 19712 24544 19718
rect 24492 19654 24544 19660
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24320 15150 24440 15178
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24412 11150 24440 15150
rect 24504 14346 24532 19654
rect 24596 17678 24624 21830
rect 24688 21593 24716 22510
rect 24674 21584 24730 21593
rect 24674 21519 24730 21528
rect 24872 20618 24900 22918
rect 25240 22778 25268 23462
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25044 22432 25096 22438
rect 25044 22374 25096 22380
rect 25056 21690 25084 22374
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 25148 21978 25176 22102
rect 25424 22098 25452 22918
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 25148 21950 25452 21978
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24872 20590 24992 20618
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24780 18766 24808 19110
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24492 13864 24544 13870
rect 24490 13832 24492 13841
rect 24544 13832 24546 13841
rect 24490 13767 24546 13776
rect 24596 12434 24624 16594
rect 24674 16552 24730 16561
rect 24674 16487 24676 16496
rect 24728 16487 24730 16496
rect 24676 16458 24728 16464
rect 24674 16144 24730 16153
rect 24674 16079 24676 16088
rect 24728 16079 24730 16088
rect 24676 16050 24728 16056
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24688 13734 24716 15098
rect 24780 15065 24808 18226
rect 24766 15056 24822 15065
rect 24766 14991 24822 15000
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24872 13394 24900 18838
rect 24964 18426 24992 20590
rect 25056 20058 25084 21490
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25056 18358 25084 18566
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24504 12406 24624 12434
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24308 9444 24360 9450
rect 24308 9386 24360 9392
rect 24044 8894 24164 8922
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24044 4622 24072 8298
rect 24136 5710 24164 8894
rect 24320 6798 24348 9386
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24412 8090 24440 8842
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24504 6322 24532 12406
rect 24688 12374 24716 12650
rect 24766 12608 24822 12617
rect 24766 12543 24822 12552
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 24674 12200 24730 12209
rect 24674 12135 24730 12144
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11354 24624 11494
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24688 10606 24716 12135
rect 24780 11694 24808 12543
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24964 11506 24992 17546
rect 25148 15994 25176 19858
rect 25240 19310 25268 20198
rect 25332 19854 25360 21830
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25240 18834 25268 19246
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25332 18698 25360 19790
rect 25424 19514 25452 21950
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25320 18692 25372 18698
rect 25320 18634 25372 18640
rect 25424 17270 25452 19450
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 25412 17060 25464 17066
rect 25412 17002 25464 17008
rect 25056 15966 25176 15994
rect 25228 15972 25280 15978
rect 25056 15162 25084 15966
rect 25228 15914 25280 15920
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 25148 15162 25176 15846
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25056 12850 25084 14350
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25148 12986 25176 13330
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 24964 11478 25084 11506
rect 24950 11384 25006 11393
rect 24950 11319 25006 11328
rect 24964 11218 24992 11319
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24582 10160 24638 10169
rect 24582 10095 24638 10104
rect 24596 8430 24624 10095
rect 24780 9518 24808 10911
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24872 10577 24900 10678
rect 24858 10568 24914 10577
rect 24858 10503 24914 10512
rect 25056 10146 25084 11478
rect 25136 10532 25188 10538
rect 25136 10474 25188 10480
rect 24872 10118 25084 10146
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24688 7342 24716 8871
rect 24872 8650 24900 10118
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24950 9344 25006 9353
rect 24950 9279 25006 9288
rect 24964 9042 24992 9279
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24872 8622 24992 8650
rect 24860 8560 24912 8566
rect 24858 8528 24860 8537
rect 24912 8528 24914 8537
rect 24858 8463 24914 8472
rect 24964 8242 24992 8622
rect 24872 8214 24992 8242
rect 24872 7818 24900 8214
rect 24950 8120 25006 8129
rect 24950 8055 25006 8064
rect 24964 7954 24992 8055
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 24688 5166 24716 6423
rect 24780 6254 24808 7647
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24872 7313 24900 7414
rect 24858 7304 24914 7313
rect 25056 7274 25084 9998
rect 25148 9926 25176 10474
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 24858 7239 24914 7248
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 24858 6896 24914 6905
rect 24858 6831 24860 6840
rect 24912 6831 24914 6840
rect 24860 6802 24912 6808
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24872 6089 24900 6326
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 24950 5672 25006 5681
rect 24950 5607 24952 5616
rect 25004 5607 25006 5616
rect 24952 5578 25004 5584
rect 24860 5296 24912 5302
rect 24766 5264 24822 5273
rect 24860 5238 24912 5244
rect 24766 5199 24822 5208
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24688 3534 24716 4422
rect 24780 4078 24808 5199
rect 24872 4865 24900 5238
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24964 4457 24992 4490
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 25056 3942 25084 6666
rect 25148 6458 25176 8842
rect 25240 8498 25268 15914
rect 25318 15464 25374 15473
rect 25318 15399 25374 15408
rect 25332 15026 25360 15399
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25424 7546 25452 17002
rect 25608 14346 25636 23530
rect 26054 21584 26110 21593
rect 26054 21519 26110 21528
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 25700 9110 25728 21286
rect 26068 9178 26096 21519
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25134 4040 25190 4049
rect 25134 3975 25190 3984
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24964 3233 24992 3402
rect 24950 3224 25006 3233
rect 24950 3159 25006 3168
rect 25148 3126 25176 3975
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 24872 2825 24900 3062
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 22190 1592 22246 1601
rect 22190 1527 22246 1536
rect 22098 1184 22154 1193
rect 22020 1142 22098 1170
rect 22098 1119 22154 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 23400 377 23428 2450
rect 24950 2408 25006 2417
rect 24950 2343 24952 2352
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 25056 785 25084 2926
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 23386 368 23442 377
rect 23386 303 23442 312
<< via2 >>
rect 938 23724 994 23760
rect 938 23704 940 23724
rect 940 23704 992 23724
rect 992 23704 994 23724
rect 938 22636 994 22672
rect 938 22616 940 22636
rect 940 22616 992 22636
rect 992 22616 994 22636
rect 2134 24928 2190 24984
rect 2778 25880 2834 25936
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 3422 24792 3478 24848
rect 3790 23024 3846 23080
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3330 18944 3386 19000
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3238 17584 3294 17640
rect 4526 24248 4582 24304
rect 4710 23160 4766 23216
rect 3974 19896 4030 19952
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 4342 22344 4398 22400
rect 4434 22208 4490 22264
rect 4710 22208 4766 22264
rect 4802 21548 4858 21584
rect 4802 21528 4804 21548
rect 4804 21528 4856 21548
rect 4856 21528 4858 21548
rect 5170 24792 5226 24848
rect 4710 18148 4766 18184
rect 4710 18128 4712 18148
rect 4712 18128 4764 18148
rect 4764 18128 4766 18148
rect 5170 20304 5226 20360
rect 5446 26152 5502 26208
rect 6734 23432 6790 23488
rect 6550 22616 6606 22672
rect 5446 19352 5502 19408
rect 5630 21936 5686 21992
rect 6182 21392 6238 21448
rect 5630 20576 5686 20632
rect 5630 19216 5686 19272
rect 5998 20848 6054 20904
rect 4894 17176 4950 17232
rect 6366 21120 6422 21176
rect 6458 20440 6514 20496
rect 7102 20168 7158 20224
rect 6918 19760 6974 19816
rect 6918 19488 6974 19544
rect 6826 18264 6882 18320
rect 6274 16496 6330 16552
rect 4526 16088 4582 16144
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 6826 17060 6882 17096
rect 6826 17040 6828 17060
rect 6828 17040 6880 17060
rect 6880 17040 6882 17060
rect 7102 19488 7158 19544
rect 7102 18672 7158 18728
rect 7470 23568 7526 23624
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7562 22480 7618 22536
rect 7102 17756 7104 17776
rect 7104 17756 7156 17776
rect 7156 17756 7158 17776
rect 7102 17720 7158 17756
rect 8574 24656 8630 24712
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7838 20984 7894 21040
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8482 22888 8538 22944
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7838 18828 7894 18864
rect 7838 18808 7840 18828
rect 7840 18808 7892 18828
rect 7892 18808 7894 18828
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8390 18400 8446 18456
rect 8390 18164 8392 18184
rect 8392 18164 8444 18184
rect 8444 18164 8446 18184
rect 8390 18128 8446 18164
rect 8390 17992 8446 18048
rect 7930 17856 7986 17912
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 9126 23704 9182 23760
rect 8942 23432 8998 23488
rect 8758 22208 8814 22264
rect 9218 20576 9274 20632
rect 8942 19488 8998 19544
rect 8850 18944 8906 19000
rect 8666 18128 8722 18184
rect 8758 17856 8814 17912
rect 8574 16224 8630 16280
rect 6918 15408 6974 15464
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 8850 17196 8906 17232
rect 8850 17176 8852 17196
rect 8852 17176 8904 17196
rect 8904 17176 8906 17196
rect 9218 20168 9274 20224
rect 9218 19080 9274 19136
rect 9126 18944 9182 19000
rect 9126 18572 9128 18592
rect 9128 18572 9180 18592
rect 9180 18572 9182 18592
rect 9126 18536 9182 18572
rect 9862 21664 9918 21720
rect 9954 20848 10010 20904
rect 9494 19080 9550 19136
rect 9586 18944 9642 19000
rect 9494 18400 9550 18456
rect 9402 17448 9458 17504
rect 9310 16224 9366 16280
rect 9126 15408 9182 15464
rect 9034 14456 9090 14512
rect 8758 14320 8814 14376
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 10046 19624 10102 19680
rect 9954 16632 10010 16688
rect 10506 21800 10562 21856
rect 10322 19760 10378 19816
rect 11242 20848 11298 20904
rect 10690 19896 10746 19952
rect 10782 18944 10838 19000
rect 11058 19352 11114 19408
rect 11058 18400 11114 18456
rect 11334 20712 11390 20768
rect 11058 16360 11114 16416
rect 12530 24248 12586 24304
rect 12438 24112 12494 24168
rect 11978 22752 12034 22808
rect 11518 21120 11574 21176
rect 12346 22208 12402 22264
rect 12254 22072 12310 22128
rect 12714 23432 12770 23488
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 13726 23568 13782 23624
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12070 21684 12126 21720
rect 12070 21664 12072 21684
rect 12072 21664 12124 21684
rect 12124 21664 12126 21684
rect 12530 21664 12586 21720
rect 12438 21020 12440 21040
rect 12440 21020 12492 21040
rect 12492 21020 12494 21040
rect 12438 20984 12494 21020
rect 12530 20712 12586 20768
rect 12806 22344 12862 22400
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13450 21528 13506 21584
rect 11334 16224 11390 16280
rect 10966 15988 10968 16008
rect 10968 15988 11020 16008
rect 11020 15988 11022 16008
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 10322 15544 10378 15600
rect 10966 15952 11022 15988
rect 10966 15156 11022 15192
rect 10966 15136 10968 15156
rect 10968 15136 11020 15156
rect 11020 15136 11022 15156
rect 10782 15020 10838 15056
rect 10782 15000 10784 15020
rect 10784 15000 10836 15020
rect 10836 15000 10838 15020
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 11886 16224 11942 16280
rect 12530 18944 12586 19000
rect 12898 20712 12954 20768
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13450 19116 13452 19136
rect 13452 19116 13504 19136
rect 13504 19116 13506 19136
rect 13450 19080 13506 19116
rect 13450 18944 13506 19000
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13818 17176 13874 17232
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13174 15136 13230 15192
rect 13174 14864 13230 14920
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13450 15000 13506 15056
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 14094 21528 14150 21584
rect 14278 22344 14334 22400
rect 14554 23840 14610 23896
rect 14278 21528 14334 21584
rect 15658 23296 15714 23352
rect 14370 19916 14426 19952
rect 14370 19896 14372 19916
rect 14372 19896 14424 19916
rect 14424 19896 14426 19916
rect 14922 20576 14978 20632
rect 14830 19352 14886 19408
rect 14738 18944 14794 19000
rect 14646 16904 14702 16960
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 14462 12552 14518 12608
rect 15198 20440 15254 20496
rect 14922 18400 14978 18456
rect 15474 21664 15530 21720
rect 15198 19624 15254 19680
rect 15014 17992 15070 18048
rect 14922 16904 14978 16960
rect 15658 22344 15714 22400
rect 15566 18128 15622 18184
rect 15566 15972 15622 16008
rect 15566 15952 15568 15972
rect 15568 15952 15620 15972
rect 15620 15952 15622 15972
rect 16118 24928 16174 24984
rect 15934 22888 15990 22944
rect 15842 15952 15898 16008
rect 15106 13368 15162 13424
rect 15842 12144 15898 12200
rect 17038 24792 17094 24848
rect 16762 23432 16818 23488
rect 16762 22616 16818 22672
rect 17314 23432 17370 23488
rect 20166 26288 20222 26344
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17590 23024 17646 23080
rect 16854 21800 16910 21856
rect 16578 20984 16634 21040
rect 16210 17856 16266 17912
rect 16210 17584 16266 17640
rect 16946 21256 17002 21312
rect 16762 20868 16818 20904
rect 16762 20848 16764 20868
rect 16764 20848 16816 20868
rect 16816 20848 16818 20868
rect 16762 20712 16818 20768
rect 16578 19896 16634 19952
rect 16670 19080 16726 19136
rect 16670 18536 16726 18592
rect 16854 20168 16910 20224
rect 16762 17992 16818 18048
rect 16486 17176 16542 17232
rect 16762 16224 16818 16280
rect 17038 19352 17094 19408
rect 17038 18944 17094 19000
rect 17314 20304 17370 20360
rect 17314 19488 17370 19544
rect 18418 23568 18474 23624
rect 17958 23296 18014 23352
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17406 19352 17462 19408
rect 17314 16632 17370 16688
rect 17222 16360 17278 16416
rect 17038 15972 17094 16008
rect 17038 15952 17040 15972
rect 17040 15952 17092 15972
rect 17092 15952 17094 15972
rect 16578 12280 16634 12336
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 17222 15952 17278 16008
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18326 20032 18382 20088
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18050 19352 18106 19408
rect 17866 19216 17922 19272
rect 18694 23296 18750 23352
rect 18694 21936 18750 21992
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17774 15680 17830 15736
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18970 24656 19026 24712
rect 19338 24248 19394 24304
rect 19246 23588 19302 23624
rect 19246 23568 19248 23588
rect 19248 23568 19300 23588
rect 19300 23568 19302 23588
rect 19246 23296 19302 23352
rect 18878 21800 18934 21856
rect 18970 19216 19026 19272
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17866 11736 17922 11792
rect 17590 11192 17646 11248
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18694 13504 18750 13560
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18050 9560 18106 9616
rect 18878 13640 18934 13696
rect 19338 22752 19394 22808
rect 20258 26152 20314 26208
rect 19890 23024 19946 23080
rect 19614 22924 19616 22944
rect 19616 22924 19668 22944
rect 19668 22924 19670 22944
rect 19430 22616 19486 22672
rect 19614 22888 19670 22924
rect 19982 22888 20038 22944
rect 19982 22772 20038 22808
rect 19982 22752 19984 22772
rect 19984 22752 20036 22772
rect 20036 22752 20038 22772
rect 19522 20712 19578 20768
rect 19430 20032 19486 20088
rect 20074 22380 20076 22400
rect 20076 22380 20128 22400
rect 20128 22380 20130 22400
rect 20074 22344 20130 22380
rect 19890 20984 19946 21040
rect 19338 18808 19394 18864
rect 19430 16788 19486 16824
rect 19430 16768 19432 16788
rect 19432 16768 19484 16788
rect 19484 16768 19486 16788
rect 19246 16360 19302 16416
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19614 17856 19670 17912
rect 19798 17856 19854 17912
rect 19798 16632 19854 16688
rect 20258 22752 20314 22808
rect 20166 19080 20222 19136
rect 20350 17212 20352 17232
rect 20352 17212 20404 17232
rect 20404 17212 20406 17232
rect 20350 17176 20406 17212
rect 20626 22208 20682 22264
rect 20718 21528 20774 21584
rect 20810 21392 20866 21448
rect 20534 20576 20590 20632
rect 21178 23160 21234 23216
rect 21178 22344 21234 22400
rect 20994 22072 21050 22128
rect 20902 20848 20958 20904
rect 20994 20712 21050 20768
rect 20626 19372 20682 19408
rect 20626 19352 20628 19372
rect 20628 19352 20680 19372
rect 20680 19352 20682 19372
rect 20074 11056 20130 11112
rect 19522 10260 19578 10296
rect 19522 10240 19524 10260
rect 19524 10240 19576 10260
rect 19576 10240 19578 10260
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 20810 18672 20866 18728
rect 20902 18284 20958 18320
rect 20902 18264 20904 18284
rect 20904 18264 20956 18284
rect 20956 18264 20958 18284
rect 20810 17176 20866 17232
rect 21178 18944 21234 19000
rect 21178 18264 21234 18320
rect 20810 15680 20866 15736
rect 20718 12416 20774 12472
rect 20718 11464 20774 11520
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 20810 11056 20866 11112
rect 20994 12416 21050 12472
rect 21914 25608 21970 25664
rect 21546 21120 21602 21176
rect 21546 18672 21602 18728
rect 21546 17040 21602 17096
rect 22006 22208 22062 22264
rect 21914 22072 21970 22128
rect 22466 26016 22522 26072
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 21914 21392 21970 21448
rect 22282 21936 22338 21992
rect 22190 20848 22246 20904
rect 21914 19216 21970 19272
rect 21270 12860 21272 12880
rect 21272 12860 21324 12880
rect 21324 12860 21326 12880
rect 21270 12824 21326 12860
rect 21086 11736 21142 11792
rect 21822 16632 21878 16688
rect 22742 22616 22798 22672
rect 22466 20440 22522 20496
rect 22650 19760 22706 19816
rect 22282 19080 22338 19136
rect 22190 17484 22192 17504
rect 22192 17484 22244 17504
rect 22244 17484 22246 17504
rect 22190 17448 22246 17484
rect 22006 16244 22062 16280
rect 22006 16224 22008 16244
rect 22008 16224 22060 16244
rect 22060 16224 22062 16244
rect 22466 16904 22522 16960
rect 21822 13912 21878 13968
rect 21546 9560 21602 9616
rect 22190 13368 22246 13424
rect 24950 26424 25006 26480
rect 23386 23976 23442 24032
rect 23294 22480 23350 22536
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23662 22380 23664 22400
rect 23664 22380 23716 22400
rect 23716 22380 23718 22400
rect 23662 22344 23718 22380
rect 23386 20748 23388 20768
rect 23388 20748 23440 20768
rect 23440 20748 23442 20768
rect 23386 20712 23442 20748
rect 23202 20476 23204 20496
rect 23204 20476 23256 20496
rect 23256 20476 23258 20496
rect 23202 20440 23258 20476
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22742 17992 22798 18048
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17876 23442 17912
rect 23386 17856 23388 17876
rect 23388 17856 23440 17876
rect 23440 17856 23442 17876
rect 23294 17720 23350 17776
rect 23386 17604 23442 17640
rect 23386 17584 23388 17604
rect 23388 17584 23440 17604
rect 23440 17584 23442 17604
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23386 17040 23442 17096
rect 23386 15952 23442 16008
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22742 13912 22798 13968
rect 22650 13640 22706 13696
rect 22650 12824 22706 12880
rect 22098 1944 22154 2000
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23018 12960 23074 13016
rect 22926 12860 22928 12880
rect 22928 12860 22980 12880
rect 22980 12860 22982 12880
rect 22926 12824 22982 12860
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23846 18828 23902 18864
rect 23846 18808 23848 18828
rect 23848 18808 23900 18828
rect 23900 18808 23902 18828
rect 24122 21936 24178 21992
rect 24766 25200 24822 25256
rect 24122 20984 24178 21040
rect 24030 20868 24086 20904
rect 24030 20848 24032 20868
rect 24032 20848 24084 20868
rect 24084 20848 24086 20868
rect 23386 14612 23442 14648
rect 23386 14592 23388 14612
rect 23388 14592 23440 14612
rect 23440 14592 23442 14612
rect 23754 14456 23810 14512
rect 23386 11600 23442 11656
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 23662 12824 23718 12880
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24674 21528 24730 21584
rect 24490 13812 24492 13832
rect 24492 13812 24544 13832
rect 24544 13812 24546 13832
rect 24490 13776 24546 13812
rect 24674 16516 24730 16552
rect 24674 16496 24676 16516
rect 24676 16496 24728 16516
rect 24728 16496 24730 16516
rect 24674 16108 24730 16144
rect 24674 16088 24676 16108
rect 24676 16088 24728 16108
rect 24728 16088 24730 16108
rect 24766 15000 24822 15056
rect 24766 12552 24822 12608
rect 24674 12144 24730 12200
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24950 11328 25006 11384
rect 24766 10920 24822 10976
rect 24582 10104 24638 10160
rect 24858 10512 24914 10568
rect 24674 8880 24730 8936
rect 24950 9288 25006 9344
rect 24858 8508 24860 8528
rect 24860 8508 24912 8528
rect 24912 8508 24914 8528
rect 24858 8472 24914 8508
rect 24950 8064 25006 8120
rect 24766 7656 24822 7712
rect 24674 6432 24730 6488
rect 24858 7248 24914 7304
rect 24858 6860 24914 6896
rect 24858 6840 24860 6860
rect 24860 6840 24912 6860
rect 24912 6840 24914 6860
rect 24858 6024 24914 6080
rect 24950 5636 25006 5672
rect 24950 5616 24952 5636
rect 24952 5616 25004 5636
rect 25004 5616 25006 5636
rect 24766 5208 24822 5264
rect 24858 4800 24914 4856
rect 24950 4392 25006 4448
rect 25318 15408 25374 15464
rect 26054 21528 26110 21584
rect 25134 3984 25190 4040
rect 24950 3576 25006 3632
rect 24950 3168 25006 3224
rect 24858 2760 24914 2816
rect 22190 1536 22246 1592
rect 22098 1128 22154 1184
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 25042 720 25098 776
rect 23386 312 23442 368
<< metal3 >>
rect 24945 26482 25011 26485
rect 26200 26482 27000 26512
rect 24945 26480 27000 26482
rect 24945 26424 24950 26480
rect 25006 26424 27000 26480
rect 24945 26422 27000 26424
rect 24945 26419 25011 26422
rect 26200 26392 27000 26422
rect 20161 26346 20227 26349
rect 5582 26344 20227 26346
rect 5582 26288 20166 26344
rect 20222 26288 20227 26344
rect 5582 26286 20227 26288
rect 5441 26210 5507 26213
rect 5582 26210 5642 26286
rect 20161 26283 20227 26286
rect 5441 26208 5642 26210
rect 5441 26152 5446 26208
rect 5502 26152 5642 26208
rect 5441 26150 5642 26152
rect 5441 26147 5507 26150
rect 6310 26148 6316 26212
rect 6380 26210 6386 26212
rect 20253 26210 20319 26213
rect 6380 26208 20319 26210
rect 6380 26152 20258 26208
rect 20314 26152 20319 26208
rect 6380 26150 20319 26152
rect 6380 26148 6386 26150
rect 20253 26147 20319 26150
rect 22461 26074 22527 26077
rect 26200 26074 27000 26104
rect 22461 26072 27000 26074
rect 22461 26016 22466 26072
rect 22522 26016 27000 26072
rect 22461 26014 27000 26016
rect 22461 26011 22527 26014
rect 26200 25984 27000 26014
rect 0 25938 800 25968
rect 2773 25938 2839 25941
rect 0 25936 2839 25938
rect 0 25880 2778 25936
rect 2834 25880 2839 25936
rect 0 25878 2839 25880
rect 0 25848 800 25878
rect 2773 25875 2839 25878
rect 21909 25666 21975 25669
rect 26200 25666 27000 25696
rect 21909 25664 27000 25666
rect 21909 25608 21914 25664
rect 21970 25608 27000 25664
rect 21909 25606 27000 25608
rect 21909 25603 21975 25606
rect 26200 25576 27000 25606
rect 24761 25258 24827 25261
rect 26200 25258 27000 25288
rect 24761 25256 27000 25258
rect 24761 25200 24766 25256
rect 24822 25200 27000 25256
rect 24761 25198 27000 25200
rect 24761 25195 24827 25198
rect 26200 25168 27000 25198
rect 2129 24986 2195 24989
rect 16113 24986 16179 24989
rect 2129 24984 16179 24986
rect 2129 24928 2134 24984
rect 2190 24928 16118 24984
rect 16174 24928 16179 24984
rect 2129 24926 16179 24928
rect 2129 24923 2195 24926
rect 16113 24923 16179 24926
rect 0 24850 800 24880
rect 3417 24850 3483 24853
rect 0 24848 3483 24850
rect 0 24792 3422 24848
rect 3478 24792 3483 24848
rect 0 24790 3483 24792
rect 0 24760 800 24790
rect 3417 24787 3483 24790
rect 5165 24850 5231 24853
rect 17033 24850 17099 24853
rect 26200 24850 27000 24880
rect 5165 24848 17099 24850
rect 5165 24792 5170 24848
rect 5226 24792 17038 24848
rect 17094 24792 17099 24848
rect 5165 24790 17099 24792
rect 5165 24787 5231 24790
rect 17033 24787 17099 24790
rect 22050 24790 27000 24850
rect 8569 24714 8635 24717
rect 18965 24714 19031 24717
rect 8569 24712 19031 24714
rect 8569 24656 8574 24712
rect 8630 24656 18970 24712
rect 19026 24656 19031 24712
rect 8569 24654 19031 24656
rect 8569 24651 8635 24654
rect 18965 24651 19031 24654
rect 14406 24516 14412 24580
rect 14476 24578 14482 24580
rect 22050 24578 22110 24790
rect 26200 24760 27000 24790
rect 14476 24518 22110 24578
rect 14476 24516 14482 24518
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 26200 24442 27000 24472
rect 24166 24382 27000 24442
rect 4521 24306 4587 24309
rect 12525 24306 12591 24309
rect 4521 24304 12591 24306
rect 4521 24248 4526 24304
rect 4582 24248 12530 24304
rect 12586 24248 12591 24304
rect 4521 24246 12591 24248
rect 4521 24243 4587 24246
rect 12525 24243 12591 24246
rect 19333 24308 19399 24309
rect 19333 24304 19380 24308
rect 19444 24306 19450 24308
rect 19333 24248 19338 24304
rect 19333 24244 19380 24248
rect 19444 24246 19490 24306
rect 19444 24244 19450 24246
rect 19333 24243 19399 24244
rect 12433 24170 12499 24173
rect 24166 24170 24226 24382
rect 26200 24352 27000 24382
rect 12433 24168 24226 24170
rect 12433 24112 12438 24168
rect 12494 24112 24226 24168
rect 12433 24110 24226 24112
rect 12433 24107 12499 24110
rect 23381 24034 23447 24037
rect 26200 24034 27000 24064
rect 23381 24032 27000 24034
rect 23381 23976 23386 24032
rect 23442 23976 27000 24032
rect 23381 23974 27000 23976
rect 23381 23971 23447 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 8518 23836 8524 23900
rect 8588 23898 8594 23900
rect 14549 23898 14615 23901
rect 8588 23896 14615 23898
rect 8588 23840 14554 23896
rect 14610 23840 14615 23896
rect 8588 23838 14615 23840
rect 8588 23836 8594 23838
rect 14549 23835 14615 23838
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 9121 23762 9187 23765
rect 15326 23762 15332 23764
rect 9121 23760 15332 23762
rect 9121 23704 9126 23760
rect 9182 23704 15332 23760
rect 9121 23702 15332 23704
rect 9121 23699 9187 23702
rect 15326 23700 15332 23702
rect 15396 23700 15402 23764
rect 7465 23626 7531 23629
rect 13721 23626 13787 23629
rect 7465 23624 13787 23626
rect 7465 23568 7470 23624
rect 7526 23568 13726 23624
rect 13782 23568 13787 23624
rect 7465 23566 13787 23568
rect 7465 23563 7531 23566
rect 13721 23563 13787 23566
rect 18413 23626 18479 23629
rect 19241 23626 19307 23629
rect 18413 23624 19307 23626
rect 18413 23568 18418 23624
rect 18474 23568 19246 23624
rect 19302 23568 19307 23624
rect 18413 23566 19307 23568
rect 18413 23563 18479 23566
rect 19241 23563 19307 23566
rect 21214 23564 21220 23628
rect 21284 23626 21290 23628
rect 26200 23626 27000 23656
rect 21284 23566 27000 23626
rect 21284 23564 21290 23566
rect 26200 23536 27000 23566
rect 6729 23492 6795 23493
rect 6678 23490 6684 23492
rect 6638 23430 6684 23490
rect 6748 23488 6795 23492
rect 6790 23432 6795 23488
rect 6678 23428 6684 23430
rect 6748 23428 6795 23432
rect 6729 23427 6795 23428
rect 8937 23490 9003 23493
rect 12709 23490 12775 23493
rect 8937 23488 12775 23490
rect 8937 23432 8942 23488
rect 8998 23432 12714 23488
rect 12770 23432 12775 23488
rect 8937 23430 12775 23432
rect 8937 23427 9003 23430
rect 12709 23427 12775 23430
rect 14590 23428 14596 23492
rect 14660 23490 14666 23492
rect 16757 23490 16823 23493
rect 14660 23488 16823 23490
rect 14660 23432 16762 23488
rect 16818 23432 16823 23488
rect 14660 23430 16823 23432
rect 14660 23428 14666 23430
rect 16757 23427 16823 23430
rect 17309 23492 17375 23493
rect 17309 23488 17356 23492
rect 17420 23490 17426 23492
rect 17309 23432 17314 23488
rect 17309 23428 17356 23432
rect 17420 23430 17466 23490
rect 17420 23428 17426 23430
rect 17309 23427 17375 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 15653 23354 15719 23357
rect 17953 23354 18019 23357
rect 18689 23354 18755 23357
rect 19241 23354 19307 23357
rect 15653 23352 19307 23354
rect 15653 23296 15658 23352
rect 15714 23296 17958 23352
rect 18014 23296 18694 23352
rect 18750 23296 19246 23352
rect 19302 23296 19307 23352
rect 15653 23294 19307 23296
rect 15653 23291 15719 23294
rect 17953 23291 18019 23294
rect 18689 23291 18755 23294
rect 19241 23291 19307 23294
rect 4705 23218 4771 23221
rect 21173 23218 21239 23221
rect 4705 23216 21239 23218
rect 4705 23160 4710 23216
rect 4766 23160 21178 23216
rect 21234 23160 21239 23216
rect 4705 23158 21239 23160
rect 4705 23155 4771 23158
rect 21173 23155 21239 23158
rect 22686 23156 22692 23220
rect 22756 23218 22762 23220
rect 26200 23218 27000 23248
rect 22756 23158 27000 23218
rect 22756 23156 22762 23158
rect 26200 23128 27000 23158
rect 3785 23082 3851 23085
rect 17585 23082 17651 23085
rect 19885 23082 19951 23085
rect 3785 23080 17651 23082
rect 3785 23024 3790 23080
rect 3846 23024 17590 23080
rect 17646 23024 17651 23080
rect 3785 23022 17651 23024
rect 3785 23019 3851 23022
rect 17585 23019 17651 23022
rect 17726 23080 19951 23082
rect 17726 23024 19890 23080
rect 19946 23024 19951 23080
rect 17726 23022 19951 23024
rect 8477 22946 8543 22949
rect 15929 22946 15995 22949
rect 8477 22944 15995 22946
rect 8477 22888 8482 22944
rect 8538 22888 15934 22944
rect 15990 22888 15995 22944
rect 8477 22886 15995 22888
rect 8477 22883 8543 22886
rect 15929 22883 15995 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 11973 22810 12039 22813
rect 17726 22810 17786 23022
rect 19885 23019 19951 23022
rect 19609 22946 19675 22949
rect 19977 22946 20043 22949
rect 19609 22944 20043 22946
rect 19609 22888 19614 22944
rect 19670 22888 19982 22944
rect 20038 22888 20043 22944
rect 19609 22886 20043 22888
rect 19609 22883 19675 22886
rect 19977 22883 20043 22886
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 11973 22808 17786 22810
rect 11973 22752 11978 22808
rect 12034 22752 17786 22808
rect 11973 22750 17786 22752
rect 19333 22810 19399 22813
rect 19977 22810 20043 22813
rect 19333 22808 20043 22810
rect 19333 22752 19338 22808
rect 19394 22752 19982 22808
rect 20038 22752 20043 22808
rect 19333 22750 20043 22752
rect 11973 22747 12039 22750
rect 19333 22747 19399 22750
rect 19977 22747 20043 22750
rect 20253 22810 20319 22813
rect 26200 22810 27000 22840
rect 20253 22808 27000 22810
rect 20253 22752 20258 22808
rect 20314 22752 27000 22808
rect 20253 22750 27000 22752
rect 20253 22747 20319 22750
rect 26200 22720 27000 22750
rect 0 22674 800 22704
rect 933 22674 999 22677
rect 0 22672 999 22674
rect 0 22616 938 22672
rect 994 22616 999 22672
rect 0 22614 999 22616
rect 0 22584 800 22614
rect 933 22611 999 22614
rect 6545 22674 6611 22677
rect 16757 22674 16823 22677
rect 6545 22672 16823 22674
rect 6545 22616 6550 22672
rect 6606 22616 16762 22672
rect 16818 22616 16823 22672
rect 6545 22614 16823 22616
rect 6545 22611 6611 22614
rect 16757 22611 16823 22614
rect 19425 22674 19491 22677
rect 22737 22674 22803 22677
rect 19425 22672 22803 22674
rect 19425 22616 19430 22672
rect 19486 22616 22742 22672
rect 22798 22616 22803 22672
rect 19425 22614 22803 22616
rect 19425 22611 19491 22614
rect 22737 22611 22803 22614
rect 7557 22538 7623 22541
rect 7557 22536 16498 22538
rect 7557 22480 7562 22536
rect 7618 22480 16498 22536
rect 7557 22478 16498 22480
rect 7557 22475 7623 22478
rect 4337 22402 4403 22405
rect 12801 22402 12867 22405
rect 4337 22400 12867 22402
rect 4337 22344 4342 22400
rect 4398 22344 12806 22400
rect 12862 22344 12867 22400
rect 4337 22342 12867 22344
rect 4337 22339 4403 22342
rect 12801 22339 12867 22342
rect 14273 22402 14339 22405
rect 15653 22402 15719 22405
rect 14273 22400 15719 22402
rect 14273 22344 14278 22400
rect 14334 22344 15658 22400
rect 15714 22344 15719 22400
rect 14273 22342 15719 22344
rect 14273 22339 14339 22342
rect 15653 22339 15719 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 4429 22266 4495 22269
rect 4705 22266 4771 22269
rect 4429 22264 4771 22266
rect 4429 22208 4434 22264
rect 4490 22208 4710 22264
rect 4766 22208 4771 22264
rect 4429 22206 4771 22208
rect 4429 22203 4495 22206
rect 4705 22203 4771 22206
rect 8753 22266 8819 22269
rect 12341 22266 12407 22269
rect 8753 22264 12407 22266
rect 8753 22208 8758 22264
rect 8814 22208 12346 22264
rect 12402 22208 12407 22264
rect 8753 22206 12407 22208
rect 16438 22266 16498 22478
rect 19190 22476 19196 22540
rect 19260 22538 19266 22540
rect 23289 22538 23355 22541
rect 19260 22536 23355 22538
rect 19260 22480 23294 22536
rect 23350 22480 23355 22536
rect 19260 22478 23355 22480
rect 19260 22476 19266 22478
rect 23289 22475 23355 22478
rect 19926 22340 19932 22404
rect 19996 22402 20002 22404
rect 20069 22402 20135 22405
rect 19996 22400 20135 22402
rect 19996 22344 20074 22400
rect 20130 22344 20135 22400
rect 19996 22342 20135 22344
rect 19996 22340 20002 22342
rect 20069 22339 20135 22342
rect 21173 22402 21239 22405
rect 23657 22404 23723 22405
rect 21173 22400 21834 22402
rect 21173 22344 21178 22400
rect 21234 22344 21834 22400
rect 21173 22342 21834 22344
rect 21173 22339 21239 22342
rect 20621 22266 20687 22269
rect 16438 22264 20687 22266
rect 16438 22208 20626 22264
rect 20682 22208 20687 22264
rect 16438 22206 20687 22208
rect 8753 22203 8819 22206
rect 12341 22203 12407 22206
rect 20621 22203 20687 22206
rect 12249 22130 12315 22133
rect 20989 22130 21055 22133
rect 12249 22128 21055 22130
rect 12249 22072 12254 22128
rect 12310 22072 20994 22128
rect 21050 22072 21055 22128
rect 12249 22070 21055 22072
rect 21774 22130 21834 22342
rect 23606 22340 23612 22404
rect 23676 22402 23723 22404
rect 26200 22402 27000 22432
rect 23676 22400 23768 22402
rect 23718 22344 23768 22400
rect 23676 22342 23768 22344
rect 24350 22342 27000 22402
rect 23676 22340 23723 22342
rect 23657 22339 23723 22340
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 22001 22268 22067 22269
rect 21950 22266 21956 22268
rect 21910 22206 21956 22266
rect 22020 22264 22067 22268
rect 22062 22208 22067 22264
rect 21950 22204 21956 22206
rect 22020 22204 22067 22208
rect 22001 22203 22067 22204
rect 21909 22130 21975 22133
rect 24350 22130 24410 22342
rect 26200 22312 27000 22342
rect 21774 22128 21975 22130
rect 21774 22072 21914 22128
rect 21970 22072 21975 22128
rect 21774 22070 21975 22072
rect 12249 22067 12315 22070
rect 20989 22067 21055 22070
rect 21909 22067 21975 22070
rect 22326 22070 24410 22130
rect 22326 21997 22386 22070
rect 5625 21994 5691 21997
rect 18689 21994 18755 21997
rect 5625 21992 18755 21994
rect 5625 21936 5630 21992
rect 5686 21936 18694 21992
rect 18750 21936 18755 21992
rect 5625 21934 18755 21936
rect 5625 21931 5691 21934
rect 18689 21931 18755 21934
rect 22277 21992 22386 21997
rect 22277 21936 22282 21992
rect 22338 21936 22386 21992
rect 22277 21934 22386 21936
rect 24117 21994 24183 21997
rect 26200 21994 27000 22024
rect 24117 21992 27000 21994
rect 24117 21936 24122 21992
rect 24178 21936 27000 21992
rect 24117 21934 27000 21936
rect 22277 21931 22343 21934
rect 24117 21931 24183 21934
rect 26200 21904 27000 21934
rect 10501 21858 10567 21861
rect 16849 21858 16915 21861
rect 10501 21856 16915 21858
rect 10501 21800 10506 21856
rect 10562 21800 16854 21856
rect 16910 21800 16915 21856
rect 10501 21798 16915 21800
rect 10501 21795 10567 21798
rect 16849 21795 16915 21798
rect 18454 21796 18460 21860
rect 18524 21858 18530 21860
rect 18873 21858 18939 21861
rect 18524 21856 18939 21858
rect 18524 21800 18878 21856
rect 18934 21800 18939 21856
rect 18524 21798 18939 21800
rect 18524 21796 18530 21798
rect 18873 21795 18939 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 9857 21722 9923 21725
rect 12065 21722 12131 21725
rect 9857 21720 12131 21722
rect 9857 21664 9862 21720
rect 9918 21664 12070 21720
rect 12126 21664 12131 21720
rect 9857 21662 12131 21664
rect 9857 21659 9923 21662
rect 12065 21659 12131 21662
rect 12525 21722 12591 21725
rect 15469 21722 15535 21725
rect 12525 21720 15535 21722
rect 12525 21664 12530 21720
rect 12586 21664 15474 21720
rect 15530 21664 15535 21720
rect 12525 21662 15535 21664
rect 12525 21659 12591 21662
rect 15469 21659 15535 21662
rect 4797 21586 4863 21589
rect 13445 21586 13511 21589
rect 4797 21584 13511 21586
rect 4797 21528 4802 21584
rect 4858 21528 13450 21584
rect 13506 21528 13511 21584
rect 4797 21526 13511 21528
rect 4797 21523 4863 21526
rect 13445 21523 13511 21526
rect 14089 21586 14155 21589
rect 14273 21586 14339 21589
rect 14089 21584 14339 21586
rect 14089 21528 14094 21584
rect 14150 21528 14278 21584
rect 14334 21528 14339 21584
rect 14089 21526 14339 21528
rect 14089 21523 14155 21526
rect 14273 21523 14339 21526
rect 20713 21586 20779 21589
rect 24669 21586 24735 21589
rect 20713 21584 24735 21586
rect 20713 21528 20718 21584
rect 20774 21528 24674 21584
rect 24730 21528 24735 21584
rect 20713 21526 24735 21528
rect 20713 21523 20779 21526
rect 24669 21523 24735 21526
rect 26049 21586 26115 21589
rect 26200 21586 27000 21616
rect 26049 21584 27000 21586
rect 26049 21528 26054 21584
rect 26110 21528 27000 21584
rect 26049 21526 27000 21528
rect 26049 21523 26115 21526
rect 26200 21496 27000 21526
rect 6177 21450 6243 21453
rect 19374 21450 19380 21452
rect 6177 21448 19380 21450
rect 6177 21392 6182 21448
rect 6238 21392 19380 21448
rect 6177 21390 19380 21392
rect 6177 21387 6243 21390
rect 19374 21388 19380 21390
rect 19444 21388 19450 21452
rect 20662 21388 20668 21452
rect 20732 21450 20738 21452
rect 20805 21450 20871 21453
rect 20732 21448 20871 21450
rect 20732 21392 20810 21448
rect 20866 21392 20871 21448
rect 20732 21390 20871 21392
rect 20732 21388 20738 21390
rect 20805 21387 20871 21390
rect 21909 21450 21975 21453
rect 21909 21448 24226 21450
rect 21909 21392 21914 21448
rect 21970 21392 24226 21448
rect 21909 21390 24226 21392
rect 21909 21387 21975 21390
rect 16430 21252 16436 21316
rect 16500 21314 16506 21316
rect 16941 21314 17007 21317
rect 16500 21312 17007 21314
rect 16500 21256 16946 21312
rect 17002 21256 17007 21312
rect 16500 21254 17007 21256
rect 16500 21252 16506 21254
rect 16941 21251 17007 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 6361 21178 6427 21181
rect 11513 21178 11579 21181
rect 21541 21178 21607 21181
rect 6361 21176 11579 21178
rect 6361 21120 6366 21176
rect 6422 21120 11518 21176
rect 11574 21120 11579 21176
rect 6361 21118 11579 21120
rect 6361 21115 6427 21118
rect 11513 21115 11579 21118
rect 13494 21176 21607 21178
rect 13494 21120 21546 21176
rect 21602 21120 21607 21176
rect 13494 21118 21607 21120
rect 24166 21178 24226 21390
rect 26200 21178 27000 21208
rect 24166 21118 27000 21178
rect 7833 21042 7899 21045
rect 12433 21042 12499 21045
rect 7833 21040 12499 21042
rect 7833 20984 7838 21040
rect 7894 20984 12438 21040
rect 12494 20984 12499 21040
rect 7833 20982 12499 20984
rect 7833 20979 7899 20982
rect 12433 20979 12499 20982
rect 12566 20980 12572 21044
rect 12636 21042 12642 21044
rect 13494 21042 13554 21118
rect 21541 21115 21607 21118
rect 26200 21088 27000 21118
rect 12636 20982 13554 21042
rect 16573 21042 16639 21045
rect 19885 21042 19951 21045
rect 24117 21042 24183 21045
rect 16573 21040 19951 21042
rect 16573 20984 16578 21040
rect 16634 20984 19890 21040
rect 19946 20984 19951 21040
rect 16573 20982 19951 20984
rect 12636 20980 12642 20982
rect 16573 20979 16639 20982
rect 19885 20979 19951 20982
rect 22326 21040 24183 21042
rect 22326 20984 24122 21040
rect 24178 20984 24183 21040
rect 22326 20982 24183 20984
rect 5993 20906 6059 20909
rect 9949 20906 10015 20909
rect 5993 20904 10015 20906
rect 5993 20848 5998 20904
rect 6054 20848 9954 20904
rect 10010 20848 10015 20904
rect 5993 20846 10015 20848
rect 5993 20843 6059 20846
rect 9949 20843 10015 20846
rect 11237 20906 11303 20909
rect 16757 20906 16823 20909
rect 20897 20906 20963 20909
rect 11237 20904 16823 20906
rect 11237 20848 11242 20904
rect 11298 20848 16762 20904
rect 16818 20848 16823 20904
rect 11237 20846 16823 20848
rect 11237 20843 11303 20846
rect 16757 20843 16823 20846
rect 16990 20904 20963 20906
rect 16990 20848 20902 20904
rect 20958 20848 20963 20904
rect 16990 20846 20963 20848
rect 11329 20770 11395 20773
rect 12382 20770 12388 20772
rect 11329 20768 12388 20770
rect 11329 20712 11334 20768
rect 11390 20712 12388 20768
rect 11329 20710 12388 20712
rect 11329 20707 11395 20710
rect 12382 20708 12388 20710
rect 12452 20708 12458 20772
rect 12525 20770 12591 20773
rect 12893 20770 12959 20773
rect 12525 20768 12959 20770
rect 12525 20712 12530 20768
rect 12586 20712 12898 20768
rect 12954 20712 12959 20768
rect 12525 20710 12959 20712
rect 12525 20707 12591 20710
rect 12893 20707 12959 20710
rect 16757 20770 16823 20773
rect 16990 20770 17050 20846
rect 20897 20843 20963 20846
rect 22185 20906 22251 20909
rect 22326 20906 22386 20982
rect 24117 20979 24183 20982
rect 22185 20904 22386 20906
rect 22185 20848 22190 20904
rect 22246 20848 22386 20904
rect 22185 20846 22386 20848
rect 22185 20843 22251 20846
rect 23422 20844 23428 20908
rect 23492 20906 23498 20908
rect 24025 20906 24091 20909
rect 23492 20904 24091 20906
rect 23492 20848 24030 20904
rect 24086 20848 24091 20904
rect 23492 20846 24091 20848
rect 23492 20844 23498 20846
rect 24025 20843 24091 20846
rect 16757 20768 17050 20770
rect 16757 20712 16762 20768
rect 16818 20712 17050 20768
rect 16757 20710 17050 20712
rect 19517 20770 19583 20773
rect 20989 20770 21055 20773
rect 19517 20768 21055 20770
rect 19517 20712 19522 20768
rect 19578 20712 20994 20768
rect 21050 20712 21055 20768
rect 19517 20710 21055 20712
rect 16757 20707 16823 20710
rect 19517 20707 19583 20710
rect 20989 20707 21055 20710
rect 23381 20770 23447 20773
rect 26200 20770 27000 20800
rect 23381 20768 27000 20770
rect 23381 20712 23386 20768
rect 23442 20712 27000 20768
rect 23381 20710 27000 20712
rect 23381 20707 23447 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 26200 20680 27000 20710
rect 17946 20639 18262 20640
rect 5625 20634 5691 20637
rect 6310 20634 6316 20636
rect 5625 20632 6316 20634
rect 5625 20576 5630 20632
rect 5686 20576 6316 20632
rect 5625 20574 6316 20576
rect 5625 20571 5691 20574
rect 6310 20572 6316 20574
rect 6380 20572 6386 20636
rect 9213 20634 9279 20637
rect 14917 20634 14983 20637
rect 9213 20632 14983 20634
rect 9213 20576 9218 20632
rect 9274 20576 14922 20632
rect 14978 20576 14983 20632
rect 9213 20574 14983 20576
rect 9213 20571 9279 20574
rect 14917 20571 14983 20574
rect 19558 20572 19564 20636
rect 19628 20634 19634 20636
rect 20529 20634 20595 20637
rect 19628 20632 20595 20634
rect 19628 20576 20534 20632
rect 20590 20576 20595 20632
rect 19628 20574 20595 20576
rect 19628 20572 19634 20574
rect 20529 20571 20595 20574
rect 6453 20498 6519 20501
rect 15193 20498 15259 20501
rect 22461 20498 22527 20501
rect 23197 20498 23263 20501
rect 6453 20496 15259 20498
rect 6453 20440 6458 20496
rect 6514 20440 15198 20496
rect 15254 20440 15259 20496
rect 6453 20438 15259 20440
rect 6453 20435 6519 20438
rect 15193 20435 15259 20438
rect 17174 20496 23263 20498
rect 17174 20440 22466 20496
rect 22522 20440 23202 20496
rect 23258 20440 23263 20496
rect 17174 20438 23263 20440
rect 5165 20362 5231 20365
rect 17174 20362 17234 20438
rect 22461 20435 22527 20438
rect 23197 20435 23263 20438
rect 5165 20360 17234 20362
rect 5165 20304 5170 20360
rect 5226 20304 17234 20360
rect 5165 20302 17234 20304
rect 17309 20362 17375 20365
rect 26200 20362 27000 20392
rect 17309 20360 27000 20362
rect 17309 20304 17314 20360
rect 17370 20304 27000 20360
rect 17309 20302 27000 20304
rect 5165 20299 5231 20302
rect 17309 20299 17375 20302
rect 26200 20272 27000 20302
rect 7097 20226 7163 20229
rect 9213 20226 9279 20229
rect 7097 20224 9279 20226
rect 7097 20168 7102 20224
rect 7158 20168 9218 20224
rect 9274 20168 9279 20224
rect 7097 20166 9279 20168
rect 7097 20163 7163 20166
rect 9213 20163 9279 20166
rect 16849 20226 16915 20229
rect 16849 20224 22754 20226
rect 16849 20168 16854 20224
rect 16910 20168 22754 20224
rect 16849 20166 22754 20168
rect 16849 20163 16915 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 15142 20028 15148 20092
rect 15212 20090 15218 20092
rect 18321 20090 18387 20093
rect 19425 20092 19491 20093
rect 19374 20090 19380 20092
rect 15212 20088 18387 20090
rect 15212 20032 18326 20088
rect 18382 20032 18387 20088
rect 15212 20030 18387 20032
rect 19334 20030 19380 20090
rect 19444 20088 19491 20092
rect 19486 20032 19491 20088
rect 15212 20028 15218 20030
rect 18321 20027 18387 20030
rect 19374 20028 19380 20030
rect 19444 20028 19491 20032
rect 19425 20027 19491 20028
rect 3969 19954 4035 19957
rect 10685 19954 10751 19957
rect 14365 19954 14431 19957
rect 3969 19952 10610 19954
rect 3969 19896 3974 19952
rect 4030 19896 10610 19952
rect 3969 19894 10610 19896
rect 3969 19891 4035 19894
rect 6913 19818 6979 19821
rect 10317 19818 10383 19821
rect 6913 19816 10383 19818
rect 6913 19760 6918 19816
rect 6974 19760 10322 19816
rect 10378 19760 10383 19816
rect 6913 19758 10383 19760
rect 10550 19818 10610 19894
rect 10685 19952 14431 19954
rect 10685 19896 10690 19952
rect 10746 19896 14370 19952
rect 14426 19896 14431 19952
rect 10685 19894 14431 19896
rect 10685 19891 10751 19894
rect 14365 19891 14431 19894
rect 16573 19954 16639 19957
rect 22694 19954 22754 20166
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 26200 19954 27000 19984
rect 16573 19952 22386 19954
rect 16573 19896 16578 19952
rect 16634 19896 22386 19952
rect 16573 19894 22386 19896
rect 22694 19894 27000 19954
rect 16573 19891 16639 19894
rect 22326 19818 22386 19894
rect 26200 19864 27000 19894
rect 22645 19818 22711 19821
rect 10550 19758 22110 19818
rect 22326 19816 22711 19818
rect 22326 19760 22650 19816
rect 22706 19760 22711 19816
rect 22326 19758 22711 19760
rect 6913 19755 6979 19758
rect 10317 19755 10383 19758
rect 10041 19682 10107 19685
rect 15193 19682 15259 19685
rect 10041 19680 15259 19682
rect 10041 19624 10046 19680
rect 10102 19624 15198 19680
rect 15254 19624 15259 19680
rect 10041 19622 15259 19624
rect 10041 19619 10107 19622
rect 15193 19619 15259 19622
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 6913 19546 6979 19549
rect 7097 19546 7163 19549
rect 6913 19544 7163 19546
rect 6913 19488 6918 19544
rect 6974 19488 7102 19544
rect 7158 19488 7163 19544
rect 6913 19486 7163 19488
rect 6913 19483 6979 19486
rect 7097 19483 7163 19486
rect 8937 19546 9003 19549
rect 17309 19546 17375 19549
rect 8937 19544 17375 19546
rect 8937 19488 8942 19544
rect 8998 19488 17314 19544
rect 17370 19488 17375 19544
rect 8937 19486 17375 19488
rect 8937 19483 9003 19486
rect 17309 19483 17375 19486
rect 5441 19410 5507 19413
rect 11053 19410 11119 19413
rect 5441 19408 11119 19410
rect 5441 19352 5446 19408
rect 5502 19352 11058 19408
rect 11114 19352 11119 19408
rect 5441 19350 11119 19352
rect 5441 19347 5507 19350
rect 11053 19347 11119 19350
rect 14825 19410 14891 19413
rect 17033 19410 17099 19413
rect 14825 19408 17099 19410
rect 14825 19352 14830 19408
rect 14886 19352 17038 19408
rect 17094 19352 17099 19408
rect 14825 19350 17099 19352
rect 14825 19347 14891 19350
rect 17033 19347 17099 19350
rect 17401 19410 17467 19413
rect 18045 19410 18111 19413
rect 20621 19410 20687 19413
rect 17401 19408 20687 19410
rect 17401 19352 17406 19408
rect 17462 19352 18050 19408
rect 18106 19352 20626 19408
rect 20682 19352 20687 19408
rect 17401 19350 20687 19352
rect 17401 19347 17467 19350
rect 18045 19347 18111 19350
rect 20621 19347 20687 19350
rect 5625 19274 5691 19277
rect 17861 19274 17927 19277
rect 5625 19272 17927 19274
rect 5625 19216 5630 19272
rect 5686 19216 17866 19272
rect 17922 19216 17927 19272
rect 5625 19214 17927 19216
rect 5625 19211 5691 19214
rect 17861 19211 17927 19214
rect 18965 19274 19031 19277
rect 21909 19274 21975 19277
rect 18965 19272 21975 19274
rect 18965 19216 18970 19272
rect 19026 19216 21914 19272
rect 21970 19216 21975 19272
rect 18965 19214 21975 19216
rect 22050 19274 22110 19758
rect 22645 19755 22711 19758
rect 22318 19484 22324 19548
rect 22388 19546 22394 19548
rect 26200 19546 27000 19576
rect 22388 19486 27000 19546
rect 22388 19484 22394 19486
rect 26200 19456 27000 19486
rect 22050 19214 23490 19274
rect 18965 19211 19031 19214
rect 21909 19211 21975 19214
rect 9213 19138 9279 19141
rect 9489 19138 9555 19141
rect 9213 19136 9555 19138
rect 9213 19080 9218 19136
rect 9274 19080 9494 19136
rect 9550 19080 9555 19136
rect 9213 19078 9555 19080
rect 9213 19075 9279 19078
rect 9489 19075 9555 19078
rect 13445 19138 13511 19141
rect 16665 19138 16731 19141
rect 20161 19138 20227 19141
rect 13445 19136 14980 19138
rect 13445 19080 13450 19136
rect 13506 19080 14980 19136
rect 13445 19078 14980 19080
rect 13445 19075 13511 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 3325 19002 3391 19005
rect 8845 19002 8911 19005
rect 3325 19000 8911 19002
rect 3325 18944 3330 19000
rect 3386 18944 8850 19000
rect 8906 18944 8911 19000
rect 3325 18942 8911 18944
rect 3325 18939 3391 18942
rect 8845 18939 8911 18942
rect 9121 19002 9187 19005
rect 9581 19002 9647 19005
rect 9121 19000 9647 19002
rect 9121 18944 9126 19000
rect 9182 18944 9586 19000
rect 9642 18944 9647 19000
rect 9121 18942 9647 18944
rect 9121 18939 9187 18942
rect 9581 18939 9647 18942
rect 10777 19002 10843 19005
rect 12525 19002 12591 19005
rect 10777 19000 12591 19002
rect 10777 18944 10782 19000
rect 10838 18944 12530 19000
rect 12586 18944 12591 19000
rect 10777 18942 12591 18944
rect 10777 18939 10843 18942
rect 12525 18939 12591 18942
rect 13445 19002 13511 19005
rect 14733 19002 14799 19005
rect 13445 19000 14799 19002
rect 13445 18944 13450 19000
rect 13506 18944 14738 19000
rect 14794 18944 14799 19000
rect 13445 18942 14799 18944
rect 14920 19002 14980 19078
rect 16665 19136 20227 19138
rect 16665 19080 16670 19136
rect 16726 19080 20166 19136
rect 20222 19080 20227 19136
rect 16665 19078 20227 19080
rect 16665 19075 16731 19078
rect 20161 19075 20227 19078
rect 21030 19076 21036 19140
rect 21100 19138 21106 19140
rect 22277 19138 22343 19141
rect 21100 19136 22343 19138
rect 21100 19080 22282 19136
rect 22338 19080 22343 19136
rect 21100 19078 22343 19080
rect 23430 19138 23490 19214
rect 26200 19138 27000 19168
rect 23430 19078 27000 19138
rect 21100 19076 21106 19078
rect 22277 19075 22343 19078
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 26200 19048 27000 19078
rect 22946 19007 23262 19008
rect 17033 19002 17099 19005
rect 21173 19002 21239 19005
rect 14920 19000 17099 19002
rect 14920 18944 17038 19000
rect 17094 18944 17099 19000
rect 14920 18942 17099 18944
rect 13445 18939 13511 18942
rect 14733 18939 14799 18942
rect 17033 18939 17099 18942
rect 17174 19000 21239 19002
rect 17174 18944 21178 19000
rect 21234 18944 21239 19000
rect 17174 18942 21239 18944
rect 7833 18866 7899 18869
rect 17174 18866 17234 18942
rect 21173 18939 21239 18942
rect 7833 18864 17234 18866
rect 7833 18808 7838 18864
rect 7894 18808 17234 18864
rect 7833 18806 17234 18808
rect 19333 18866 19399 18869
rect 23841 18866 23907 18869
rect 19333 18864 23907 18866
rect 19333 18808 19338 18864
rect 19394 18808 23846 18864
rect 23902 18808 23907 18864
rect 19333 18806 23907 18808
rect 7833 18803 7899 18806
rect 19333 18803 19399 18806
rect 23841 18803 23907 18806
rect 7097 18730 7163 18733
rect 20805 18730 20871 18733
rect 7097 18728 20871 18730
rect 7097 18672 7102 18728
rect 7158 18672 20810 18728
rect 20866 18672 20871 18728
rect 7097 18670 20871 18672
rect 7097 18667 7163 18670
rect 20805 18667 20871 18670
rect 21541 18730 21607 18733
rect 26200 18730 27000 18760
rect 21541 18728 27000 18730
rect 21541 18672 21546 18728
rect 21602 18672 27000 18728
rect 21541 18670 27000 18672
rect 21541 18667 21607 18670
rect 26200 18640 27000 18670
rect 9121 18594 9187 18597
rect 16665 18594 16731 18597
rect 9121 18592 16731 18594
rect 9121 18536 9126 18592
rect 9182 18536 16670 18592
rect 16726 18536 16731 18592
rect 9121 18534 16731 18536
rect 9121 18531 9187 18534
rect 16665 18531 16731 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 8385 18458 8451 18461
rect 9489 18458 9555 18461
rect 8385 18456 9555 18458
rect 8385 18400 8390 18456
rect 8446 18400 9494 18456
rect 9550 18400 9555 18456
rect 8385 18398 9555 18400
rect 8385 18395 8451 18398
rect 9489 18395 9555 18398
rect 11053 18458 11119 18461
rect 14917 18458 14983 18461
rect 11053 18456 14983 18458
rect 11053 18400 11058 18456
rect 11114 18400 14922 18456
rect 14978 18400 14983 18456
rect 11053 18398 14983 18400
rect 11053 18395 11119 18398
rect 14917 18395 14983 18398
rect 6821 18322 6887 18325
rect 20897 18322 20963 18325
rect 6821 18320 20963 18322
rect 6821 18264 6826 18320
rect 6882 18264 20902 18320
rect 20958 18264 20963 18320
rect 6821 18262 20963 18264
rect 6821 18259 6887 18262
rect 20897 18259 20963 18262
rect 21173 18322 21239 18325
rect 26200 18322 27000 18352
rect 21173 18320 27000 18322
rect 21173 18264 21178 18320
rect 21234 18264 27000 18320
rect 21173 18262 27000 18264
rect 21173 18259 21239 18262
rect 26200 18232 27000 18262
rect 4705 18186 4771 18189
rect 8385 18186 8451 18189
rect 4705 18184 8451 18186
rect 4705 18128 4710 18184
rect 4766 18128 8390 18184
rect 8446 18128 8451 18184
rect 4705 18126 8451 18128
rect 4705 18123 4771 18126
rect 8385 18123 8451 18126
rect 8661 18186 8727 18189
rect 15561 18186 15627 18189
rect 8661 18184 15627 18186
rect 8661 18128 8666 18184
rect 8722 18128 15566 18184
rect 15622 18128 15627 18184
rect 8661 18126 15627 18128
rect 8661 18123 8727 18126
rect 15561 18123 15627 18126
rect 8385 18050 8451 18053
rect 8518 18050 8524 18052
rect 8385 18048 8524 18050
rect 8385 17992 8390 18048
rect 8446 17992 8524 18048
rect 8385 17990 8524 17992
rect 8385 17987 8451 17990
rect 8518 17988 8524 17990
rect 8588 17988 8594 18052
rect 15009 18050 15075 18053
rect 16757 18050 16823 18053
rect 15009 18048 16823 18050
rect 15009 17992 15014 18048
rect 15070 17992 16762 18048
rect 16818 17992 16823 18048
rect 15009 17990 16823 17992
rect 15009 17987 15075 17990
rect 16757 17987 16823 17990
rect 22502 17988 22508 18052
rect 22572 18050 22578 18052
rect 22737 18050 22803 18053
rect 22572 18048 22803 18050
rect 22572 17992 22742 18048
rect 22798 17992 22803 18048
rect 22572 17990 22803 17992
rect 22572 17988 22578 17990
rect 22737 17987 22803 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 7925 17914 7991 17917
rect 8753 17914 8819 17917
rect 7925 17912 8819 17914
rect 7925 17856 7930 17912
rect 7986 17856 8758 17912
rect 8814 17856 8819 17912
rect 7925 17854 8819 17856
rect 7925 17851 7991 17854
rect 8753 17851 8819 17854
rect 16205 17914 16271 17917
rect 19609 17914 19675 17917
rect 16205 17912 19675 17914
rect 16205 17856 16210 17912
rect 16266 17856 19614 17912
rect 19670 17856 19675 17912
rect 16205 17854 19675 17856
rect 16205 17851 16271 17854
rect 19609 17851 19675 17854
rect 19793 17914 19859 17917
rect 20662 17914 20668 17916
rect 19793 17912 20668 17914
rect 19793 17856 19798 17912
rect 19854 17856 20668 17912
rect 19793 17854 20668 17856
rect 19793 17851 19859 17854
rect 20662 17852 20668 17854
rect 20732 17852 20738 17916
rect 23381 17914 23447 17917
rect 26200 17914 27000 17944
rect 23381 17912 27000 17914
rect 23381 17856 23386 17912
rect 23442 17856 27000 17912
rect 23381 17854 27000 17856
rect 23381 17851 23447 17854
rect 26200 17824 27000 17854
rect 7097 17778 7163 17781
rect 23289 17778 23355 17781
rect 7097 17776 23355 17778
rect 7097 17720 7102 17776
rect 7158 17720 23294 17776
rect 23350 17720 23355 17776
rect 7097 17718 23355 17720
rect 7097 17715 7163 17718
rect 23289 17715 23355 17718
rect 3233 17642 3299 17645
rect 16205 17642 16271 17645
rect 23381 17642 23447 17645
rect 3233 17640 16271 17642
rect 3233 17584 3238 17640
rect 3294 17584 16210 17640
rect 16266 17584 16271 17640
rect 3233 17582 16271 17584
rect 3233 17579 3299 17582
rect 16205 17579 16271 17582
rect 17174 17640 23447 17642
rect 17174 17584 23386 17640
rect 23442 17584 23447 17640
rect 17174 17582 23447 17584
rect 9397 17506 9463 17509
rect 17174 17506 17234 17582
rect 23381 17579 23447 17582
rect 9397 17504 17234 17506
rect 9397 17448 9402 17504
rect 9458 17448 17234 17504
rect 9397 17446 17234 17448
rect 22185 17506 22251 17509
rect 26200 17506 27000 17536
rect 22185 17504 27000 17506
rect 22185 17448 22190 17504
rect 22246 17448 27000 17504
rect 22185 17446 27000 17448
rect 9397 17443 9463 17446
rect 22185 17443 22251 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 26200 17416 27000 17446
rect 17946 17375 18262 17376
rect 15142 17370 15148 17372
rect 8342 17310 15148 17370
rect 4889 17234 4955 17237
rect 8342 17234 8402 17310
rect 15142 17308 15148 17310
rect 15212 17308 15218 17372
rect 4889 17232 8402 17234
rect 4889 17176 4894 17232
rect 4950 17176 8402 17232
rect 4889 17174 8402 17176
rect 8845 17234 8911 17237
rect 13813 17234 13879 17237
rect 16481 17234 16547 17237
rect 8845 17232 13738 17234
rect 8845 17176 8850 17232
rect 8906 17176 13738 17232
rect 8845 17174 13738 17176
rect 4889 17171 4955 17174
rect 8845 17171 8911 17174
rect 6821 17098 6887 17101
rect 13678 17098 13738 17174
rect 13813 17232 16547 17234
rect 13813 17176 13818 17232
rect 13874 17176 16486 17232
rect 16542 17176 16547 17232
rect 13813 17174 16547 17176
rect 13813 17171 13879 17174
rect 16481 17171 16547 17174
rect 20345 17234 20411 17237
rect 20805 17234 20871 17237
rect 20345 17232 20871 17234
rect 20345 17176 20350 17232
rect 20406 17176 20810 17232
rect 20866 17176 20871 17232
rect 20345 17174 20871 17176
rect 20345 17171 20411 17174
rect 20805 17171 20871 17174
rect 21541 17098 21607 17101
rect 6821 17096 13554 17098
rect 6821 17040 6826 17096
rect 6882 17040 13554 17096
rect 6821 17038 13554 17040
rect 13678 17096 21607 17098
rect 13678 17040 21546 17096
rect 21602 17040 21607 17096
rect 13678 17038 21607 17040
rect 6821 17035 6887 17038
rect 13494 16962 13554 17038
rect 21541 17035 21607 17038
rect 23381 17098 23447 17101
rect 26200 17098 27000 17128
rect 23381 17096 27000 17098
rect 23381 17040 23386 17096
rect 23442 17040 27000 17096
rect 23381 17038 27000 17040
rect 23381 17035 23447 17038
rect 26200 17008 27000 17038
rect 14641 16962 14707 16965
rect 13494 16960 14707 16962
rect 13494 16904 14646 16960
rect 14702 16904 14707 16960
rect 13494 16902 14707 16904
rect 14641 16899 14707 16902
rect 14917 16962 14983 16965
rect 22461 16962 22527 16965
rect 14917 16960 22527 16962
rect 14917 16904 14922 16960
rect 14978 16904 22466 16960
rect 22522 16904 22527 16960
rect 14917 16902 22527 16904
rect 14917 16899 14983 16902
rect 22461 16899 22527 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 15326 16764 15332 16828
rect 15396 16826 15402 16828
rect 19425 16826 19491 16829
rect 15396 16766 19258 16826
rect 15396 16764 15402 16766
rect 9949 16690 10015 16693
rect 17309 16690 17375 16693
rect 9949 16688 17375 16690
rect 9949 16632 9954 16688
rect 10010 16632 17314 16688
rect 17370 16632 17375 16688
rect 9949 16630 17375 16632
rect 19198 16690 19258 16766
rect 19425 16824 22110 16826
rect 19425 16768 19430 16824
rect 19486 16768 22110 16824
rect 19425 16766 22110 16768
rect 19425 16763 19491 16766
rect 19793 16690 19859 16693
rect 19198 16688 19859 16690
rect 19198 16632 19798 16688
rect 19854 16632 19859 16688
rect 19198 16630 19859 16632
rect 9949 16627 10015 16630
rect 17309 16627 17375 16630
rect 19793 16627 19859 16630
rect 21582 16628 21588 16692
rect 21652 16690 21658 16692
rect 21817 16690 21883 16693
rect 21652 16688 21883 16690
rect 21652 16632 21822 16688
rect 21878 16632 21883 16688
rect 21652 16630 21883 16632
rect 22050 16690 22110 16766
rect 26200 16690 27000 16720
rect 22050 16630 27000 16690
rect 21652 16628 21658 16630
rect 21817 16627 21883 16630
rect 26200 16600 27000 16630
rect 6269 16554 6335 16557
rect 24669 16554 24735 16557
rect 6269 16552 24735 16554
rect 6269 16496 6274 16552
rect 6330 16496 24674 16552
rect 24730 16496 24735 16552
rect 6269 16494 24735 16496
rect 6269 16491 6335 16494
rect 24669 16491 24735 16494
rect 11053 16418 11119 16421
rect 17217 16418 17283 16421
rect 11053 16416 17283 16418
rect 11053 16360 11058 16416
rect 11114 16360 17222 16416
rect 17278 16360 17283 16416
rect 11053 16358 17283 16360
rect 11053 16355 11119 16358
rect 17217 16355 17283 16358
rect 19241 16418 19307 16421
rect 19241 16416 24226 16418
rect 19241 16360 19246 16416
rect 19302 16360 24226 16416
rect 19241 16358 24226 16360
rect 19241 16355 19307 16358
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 8569 16282 8635 16285
rect 9305 16282 9371 16285
rect 11329 16282 11395 16285
rect 8569 16280 11395 16282
rect 8569 16224 8574 16280
rect 8630 16224 9310 16280
rect 9366 16224 11334 16280
rect 11390 16224 11395 16280
rect 8569 16222 11395 16224
rect 8569 16219 8635 16222
rect 9305 16219 9371 16222
rect 11329 16219 11395 16222
rect 11881 16282 11947 16285
rect 16757 16282 16823 16285
rect 22001 16284 22067 16285
rect 21950 16282 21956 16284
rect 11881 16280 16823 16282
rect 11881 16224 11886 16280
rect 11942 16224 16762 16280
rect 16818 16224 16823 16280
rect 11881 16222 16823 16224
rect 21910 16222 21956 16282
rect 22020 16280 22067 16284
rect 22062 16224 22067 16280
rect 11881 16219 11947 16222
rect 16757 16219 16823 16222
rect 21950 16220 21956 16222
rect 22020 16220 22067 16224
rect 24166 16282 24226 16358
rect 26200 16282 27000 16312
rect 24166 16222 27000 16282
rect 22001 16219 22067 16220
rect 26200 16192 27000 16222
rect 4521 16146 4587 16149
rect 24669 16146 24735 16149
rect 4521 16144 24735 16146
rect 4521 16088 4526 16144
rect 4582 16088 24674 16144
rect 24730 16088 24735 16144
rect 4521 16086 24735 16088
rect 4521 16083 4587 16086
rect 24669 16083 24735 16086
rect 10961 16010 11027 16013
rect 15561 16010 15627 16013
rect 10961 16008 15627 16010
rect 10961 15952 10966 16008
rect 11022 15952 15566 16008
rect 15622 15952 15627 16008
rect 10961 15950 15627 15952
rect 10961 15947 11027 15950
rect 15561 15947 15627 15950
rect 15837 16010 15903 16013
rect 17033 16010 17099 16013
rect 15837 16008 17099 16010
rect 15837 15952 15842 16008
rect 15898 15952 17038 16008
rect 17094 15952 17099 16008
rect 15837 15950 17099 15952
rect 15837 15947 15903 15950
rect 17033 15947 17099 15950
rect 17217 16010 17283 16013
rect 23381 16010 23447 16013
rect 17217 16008 23447 16010
rect 17217 15952 17222 16008
rect 17278 15952 23386 16008
rect 23442 15952 23447 16008
rect 17217 15950 23447 15952
rect 17217 15947 17283 15950
rect 23381 15947 23447 15950
rect 26200 15874 27000 15904
rect 24166 15814 27000 15874
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 17769 15738 17835 15741
rect 20805 15738 20871 15741
rect 17769 15736 20871 15738
rect 17769 15680 17774 15736
rect 17830 15680 20810 15736
rect 20866 15680 20871 15736
rect 17769 15678 20871 15680
rect 17769 15675 17835 15678
rect 20805 15675 20871 15678
rect 10317 15602 10383 15605
rect 22502 15602 22508 15604
rect 10317 15600 22508 15602
rect 10317 15544 10322 15600
rect 10378 15544 22508 15600
rect 10317 15542 22508 15544
rect 10317 15539 10383 15542
rect 22502 15540 22508 15542
rect 22572 15540 22578 15604
rect 6913 15466 6979 15469
rect 9121 15466 9187 15469
rect 16430 15466 16436 15468
rect 6913 15464 8402 15466
rect 6913 15408 6918 15464
rect 6974 15408 8402 15464
rect 6913 15406 8402 15408
rect 6913 15403 6979 15406
rect 8342 15330 8402 15406
rect 9121 15464 16436 15466
rect 9121 15408 9126 15464
rect 9182 15408 16436 15464
rect 9121 15406 16436 15408
rect 9121 15403 9187 15406
rect 16430 15404 16436 15406
rect 16500 15404 16506 15468
rect 24166 15466 24226 15814
rect 26200 15784 27000 15814
rect 17174 15406 24226 15466
rect 25313 15466 25379 15469
rect 26200 15466 27000 15496
rect 25313 15464 27000 15466
rect 25313 15408 25318 15464
rect 25374 15408 27000 15464
rect 25313 15406 27000 15408
rect 17174 15330 17234 15406
rect 25313 15403 25379 15406
rect 26200 15376 27000 15406
rect 8342 15270 17234 15330
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 10961 15194 11027 15197
rect 13169 15194 13235 15197
rect 14406 15194 14412 15196
rect 10961 15192 13235 15194
rect 10961 15136 10966 15192
rect 11022 15136 13174 15192
rect 13230 15136 13235 15192
rect 10961 15134 13235 15136
rect 10961 15131 11027 15134
rect 13169 15131 13235 15134
rect 13310 15134 14412 15194
rect 10777 15058 10843 15061
rect 13310 15058 13370 15134
rect 14406 15132 14412 15134
rect 14476 15132 14482 15196
rect 10777 15056 13370 15058
rect 10777 15000 10782 15056
rect 10838 15000 13370 15056
rect 10777 14998 13370 15000
rect 13445 15058 13511 15061
rect 23422 15058 23428 15060
rect 13445 15056 23428 15058
rect 13445 15000 13450 15056
rect 13506 15000 23428 15056
rect 13445 14998 23428 15000
rect 10777 14995 10843 14998
rect 13445 14995 13511 14998
rect 23422 14996 23428 14998
rect 23492 14996 23498 15060
rect 24761 15058 24827 15061
rect 26200 15058 27000 15088
rect 24761 15056 27000 15058
rect 24761 15000 24766 15056
rect 24822 15000 27000 15056
rect 24761 14998 27000 15000
rect 24761 14995 24827 14998
rect 26200 14968 27000 14998
rect 13169 14922 13235 14925
rect 14590 14922 14596 14924
rect 13169 14920 14596 14922
rect 13169 14864 13174 14920
rect 13230 14864 14596 14920
rect 13169 14862 14596 14864
rect 13169 14859 13235 14862
rect 14590 14860 14596 14862
rect 14660 14860 14666 14924
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 23381 14650 23447 14653
rect 26200 14650 27000 14680
rect 23381 14648 27000 14650
rect 23381 14592 23386 14648
rect 23442 14592 27000 14648
rect 23381 14590 27000 14592
rect 23381 14587 23447 14590
rect 26200 14560 27000 14590
rect 9029 14514 9095 14517
rect 23749 14514 23815 14517
rect 9029 14512 23815 14514
rect 9029 14456 9034 14512
rect 9090 14456 23754 14512
rect 23810 14456 23815 14512
rect 9029 14454 23815 14456
rect 9029 14451 9095 14454
rect 23749 14451 23815 14454
rect 8753 14378 8819 14381
rect 18454 14378 18460 14380
rect 8753 14376 18460 14378
rect 8753 14320 8758 14376
rect 8814 14320 18460 14376
rect 8753 14318 18460 14320
rect 8753 14315 8819 14318
rect 18454 14316 18460 14318
rect 18524 14316 18530 14380
rect 26200 14242 27000 14272
rect 22050 14182 27000 14242
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 21817 13970 21883 13973
rect 22050 13970 22110 14182
rect 26200 14152 27000 14182
rect 21817 13968 22110 13970
rect 21817 13912 21822 13968
rect 21878 13912 22110 13968
rect 21817 13910 22110 13912
rect 22737 13970 22803 13973
rect 22737 13968 24732 13970
rect 22737 13912 22742 13968
rect 22798 13912 24732 13968
rect 22737 13910 24732 13912
rect 21817 13907 21883 13910
rect 22737 13907 22803 13910
rect 6678 13772 6684 13836
rect 6748 13834 6754 13836
rect 24485 13834 24551 13837
rect 6748 13832 24551 13834
rect 6748 13776 24490 13832
rect 24546 13776 24551 13832
rect 6748 13774 24551 13776
rect 24672 13834 24732 13910
rect 26200 13834 27000 13864
rect 24672 13774 27000 13834
rect 6748 13772 6754 13774
rect 24485 13771 24551 13774
rect 26200 13744 27000 13774
rect 18873 13698 18939 13701
rect 22645 13698 22711 13701
rect 18873 13696 22711 13698
rect 18873 13640 18878 13696
rect 18934 13640 22650 13696
rect 22706 13640 22711 13696
rect 18873 13638 22711 13640
rect 18873 13635 18939 13638
rect 22645 13635 22711 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 18689 13562 18755 13565
rect 19190 13562 19196 13564
rect 18689 13560 19196 13562
rect 18689 13504 18694 13560
rect 18750 13504 19196 13560
rect 18689 13502 19196 13504
rect 18689 13499 18755 13502
rect 19190 13500 19196 13502
rect 19260 13500 19266 13564
rect 15101 13426 15167 13429
rect 19374 13426 19380 13428
rect 15101 13424 19380 13426
rect 15101 13368 15106 13424
rect 15162 13368 19380 13424
rect 15101 13366 19380 13368
rect 15101 13363 15167 13366
rect 19374 13364 19380 13366
rect 19444 13364 19450 13428
rect 22185 13426 22251 13429
rect 26200 13426 27000 13456
rect 22185 13424 27000 13426
rect 22185 13368 22190 13424
rect 22246 13368 27000 13424
rect 22185 13366 27000 13368
rect 22185 13363 22251 13366
rect 26200 13336 27000 13366
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 23013 13018 23079 13021
rect 26200 13018 27000 13048
rect 23013 13016 27000 13018
rect 23013 12960 23018 13016
rect 23074 12960 27000 13016
rect 23013 12958 27000 12960
rect 23013 12955 23079 12958
rect 26200 12928 27000 12958
rect 21265 12882 21331 12885
rect 22645 12882 22711 12885
rect 22921 12882 22987 12885
rect 23657 12882 23723 12885
rect 21265 12880 23723 12882
rect 21265 12824 21270 12880
rect 21326 12824 22650 12880
rect 22706 12824 22926 12880
rect 22982 12824 23662 12880
rect 23718 12824 23723 12880
rect 21265 12822 23723 12824
rect 21265 12819 21331 12822
rect 22645 12819 22711 12822
rect 22921 12819 22987 12822
rect 23657 12819 23723 12822
rect 14457 12610 14523 12613
rect 19558 12610 19564 12612
rect 14457 12608 19564 12610
rect 14457 12552 14462 12608
rect 14518 12552 19564 12608
rect 14457 12550 19564 12552
rect 14457 12547 14523 12550
rect 19558 12548 19564 12550
rect 19628 12548 19634 12612
rect 24761 12610 24827 12613
rect 26200 12610 27000 12640
rect 24761 12608 27000 12610
rect 24761 12552 24766 12608
rect 24822 12552 27000 12608
rect 24761 12550 27000 12552
rect 24761 12547 24827 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 20713 12474 20779 12477
rect 20989 12474 21055 12477
rect 20713 12472 21055 12474
rect 20713 12416 20718 12472
rect 20774 12416 20994 12472
rect 21050 12416 21055 12472
rect 20713 12414 21055 12416
rect 20713 12411 20779 12414
rect 20989 12411 21055 12414
rect 16573 12338 16639 12341
rect 21214 12338 21220 12340
rect 16573 12336 21220 12338
rect 16573 12280 16578 12336
rect 16634 12280 21220 12336
rect 16573 12278 21220 12280
rect 16573 12275 16639 12278
rect 21214 12276 21220 12278
rect 21284 12276 21290 12340
rect 15837 12202 15903 12205
rect 22686 12202 22692 12204
rect 15837 12200 22692 12202
rect 15837 12144 15842 12200
rect 15898 12144 22692 12200
rect 15837 12142 22692 12144
rect 15837 12139 15903 12142
rect 22686 12140 22692 12142
rect 22756 12140 22762 12204
rect 24669 12202 24735 12205
rect 26200 12202 27000 12232
rect 24669 12200 27000 12202
rect 24669 12144 24674 12200
rect 24730 12144 27000 12200
rect 24669 12142 27000 12144
rect 24669 12139 24735 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 20662 11868 20668 11932
rect 20732 11930 20738 11932
rect 23606 11930 23612 11932
rect 20732 11870 23612 11930
rect 20732 11868 20738 11870
rect 23606 11868 23612 11870
rect 23676 11868 23682 11932
rect 17861 11794 17927 11797
rect 21081 11794 21147 11797
rect 17861 11792 21147 11794
rect 17861 11736 17866 11792
rect 17922 11736 21086 11792
rect 21142 11736 21147 11792
rect 17861 11734 21147 11736
rect 17861 11731 17927 11734
rect 21081 11731 21147 11734
rect 24853 11794 24919 11797
rect 26200 11794 27000 11824
rect 24853 11792 27000 11794
rect 24853 11736 24858 11792
rect 24914 11736 27000 11792
rect 24853 11734 27000 11736
rect 24853 11731 24919 11734
rect 26200 11704 27000 11734
rect 23381 11658 23447 11661
rect 22694 11656 23447 11658
rect 22694 11600 23386 11656
rect 23442 11600 23447 11656
rect 22694 11598 23447 11600
rect 20713 11522 20779 11525
rect 22694 11522 22754 11598
rect 23381 11595 23447 11598
rect 20713 11520 22754 11522
rect 20713 11464 20718 11520
rect 20774 11464 22754 11520
rect 20713 11462 22754 11464
rect 20713 11459 20779 11462
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24945 11386 25011 11389
rect 26200 11386 27000 11416
rect 24945 11384 27000 11386
rect 24945 11328 24950 11384
rect 25006 11328 27000 11384
rect 24945 11326 27000 11328
rect 24945 11323 25011 11326
rect 26200 11296 27000 11326
rect 17585 11250 17651 11253
rect 22502 11250 22508 11252
rect 17585 11248 22508 11250
rect 17585 11192 17590 11248
rect 17646 11192 22508 11248
rect 17585 11190 22508 11192
rect 17585 11187 17651 11190
rect 22502 11188 22508 11190
rect 22572 11188 22578 11252
rect 19926 11052 19932 11116
rect 19996 11114 20002 11116
rect 20069 11114 20135 11117
rect 19996 11112 20135 11114
rect 19996 11056 20074 11112
rect 20130 11056 20135 11112
rect 19996 11054 20135 11056
rect 19996 11052 20002 11054
rect 20069 11051 20135 11054
rect 20805 11114 20871 11117
rect 21030 11114 21036 11116
rect 20805 11112 21036 11114
rect 20805 11056 20810 11112
rect 20866 11056 21036 11112
rect 20805 11054 21036 11056
rect 20805 11051 20871 11054
rect 21030 11052 21036 11054
rect 21100 11052 21106 11116
rect 24761 10978 24827 10981
rect 26200 10978 27000 11008
rect 24761 10976 27000 10978
rect 24761 10920 24766 10976
rect 24822 10920 27000 10976
rect 24761 10918 27000 10920
rect 24761 10915 24827 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 26200 10888 27000 10918
rect 17946 10847 18262 10848
rect 24853 10570 24919 10573
rect 26200 10570 27000 10600
rect 24853 10568 27000 10570
rect 24853 10512 24858 10568
rect 24914 10512 27000 10568
rect 24853 10510 27000 10512
rect 24853 10507 24919 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 17350 10236 17356 10300
rect 17420 10298 17426 10300
rect 19517 10298 19583 10301
rect 17420 10296 19583 10298
rect 17420 10240 19522 10296
rect 19578 10240 19583 10296
rect 17420 10238 19583 10240
rect 17420 10236 17426 10238
rect 19517 10235 19583 10238
rect 24577 10162 24643 10165
rect 26200 10162 27000 10192
rect 24577 10160 27000 10162
rect 24577 10104 24582 10160
rect 24638 10104 27000 10160
rect 24577 10102 27000 10104
rect 24577 10099 24643 10102
rect 26200 10072 27000 10102
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 18045 9618 18111 9621
rect 21541 9620 21607 9621
rect 20662 9618 20668 9620
rect 18045 9616 20668 9618
rect 18045 9560 18050 9616
rect 18106 9560 20668 9616
rect 18045 9558 20668 9560
rect 18045 9555 18111 9558
rect 20662 9556 20668 9558
rect 20732 9556 20738 9620
rect 21541 9616 21588 9620
rect 21652 9618 21658 9620
rect 21541 9560 21546 9616
rect 21541 9556 21588 9560
rect 21652 9558 21698 9618
rect 21652 9556 21658 9558
rect 21541 9555 21607 9556
rect 24945 9346 25011 9349
rect 26200 9346 27000 9376
rect 24945 9344 27000 9346
rect 24945 9288 24950 9344
rect 25006 9288 27000 9344
rect 24945 9286 27000 9288
rect 24945 9283 25011 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 24669 8938 24735 8941
rect 26200 8938 27000 8968
rect 24669 8936 27000 8938
rect 24669 8880 24674 8936
rect 24730 8880 27000 8936
rect 24669 8878 27000 8880
rect 24669 8875 24735 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24853 8530 24919 8533
rect 26200 8530 27000 8560
rect 24853 8528 27000 8530
rect 24853 8472 24858 8528
rect 24914 8472 27000 8528
rect 24853 8470 27000 8472
rect 24853 8467 24919 8470
rect 26200 8440 27000 8470
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24945 8122 25011 8125
rect 26200 8122 27000 8152
rect 24945 8120 27000 8122
rect 24945 8064 24950 8120
rect 25006 8064 27000 8120
rect 24945 8062 27000 8064
rect 24945 8059 25011 8062
rect 26200 8032 27000 8062
rect 24761 7714 24827 7717
rect 26200 7714 27000 7744
rect 24761 7712 27000 7714
rect 24761 7656 24766 7712
rect 24822 7656 27000 7712
rect 24761 7654 27000 7656
rect 24761 7651 24827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 24853 6898 24919 6901
rect 26200 6898 27000 6928
rect 24853 6896 27000 6898
rect 24853 6840 24858 6896
rect 24914 6840 27000 6896
rect 24853 6838 27000 6840
rect 24853 6835 24919 6838
rect 26200 6808 27000 6838
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 24669 6490 24735 6493
rect 26200 6490 27000 6520
rect 24669 6488 27000 6490
rect 24669 6432 24674 6488
rect 24730 6432 27000 6488
rect 24669 6430 27000 6432
rect 24669 6427 24735 6430
rect 26200 6400 27000 6430
rect 24853 6082 24919 6085
rect 26200 6082 27000 6112
rect 24853 6080 27000 6082
rect 24853 6024 24858 6080
rect 24914 6024 27000 6080
rect 24853 6022 27000 6024
rect 24853 6019 24919 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 24761 5266 24827 5269
rect 26200 5266 27000 5296
rect 24761 5264 27000 5266
rect 24761 5208 24766 5264
rect 24822 5208 27000 5264
rect 24761 5206 27000 5208
rect 24761 5203 24827 5206
rect 26200 5176 27000 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24853 4858 24919 4861
rect 26200 4858 27000 4888
rect 24853 4856 27000 4858
rect 24853 4800 24858 4856
rect 24914 4800 27000 4856
rect 24853 4798 27000 4800
rect 24853 4795 24919 4798
rect 26200 4768 27000 4798
rect 24945 4450 25011 4453
rect 26200 4450 27000 4480
rect 24945 4448 27000 4450
rect 24945 4392 24950 4448
rect 25006 4392 27000 4448
rect 24945 4390 27000 4392
rect 24945 4387 25011 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 25129 4042 25195 4045
rect 26200 4042 27000 4072
rect 25129 4040 27000 4042
rect 25129 3984 25134 4040
rect 25190 3984 27000 4040
rect 25129 3982 27000 3984
rect 25129 3979 25195 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 24945 3226 25011 3229
rect 26200 3226 27000 3256
rect 24945 3224 27000 3226
rect 24945 3168 24950 3224
rect 25006 3168 27000 3224
rect 24945 3166 27000 3168
rect 24945 3163 25011 3166
rect 26200 3136 27000 3166
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22093 2002 22159 2005
rect 26200 2002 27000 2032
rect 22093 2000 27000 2002
rect 22093 1944 22098 2000
rect 22154 1944 27000 2000
rect 22093 1942 27000 1944
rect 22093 1939 22159 1942
rect 26200 1912 27000 1942
rect 22185 1594 22251 1597
rect 26200 1594 27000 1624
rect 22185 1592 27000 1594
rect 22185 1536 22190 1592
rect 22246 1536 27000 1592
rect 22185 1534 27000 1536
rect 22185 1531 22251 1534
rect 26200 1504 27000 1534
rect 22093 1186 22159 1189
rect 26200 1186 27000 1216
rect 22093 1184 27000 1186
rect 22093 1128 22098 1184
rect 22154 1128 27000 1184
rect 22093 1126 27000 1128
rect 22093 1123 22159 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 23381 370 23447 373
rect 26200 370 27000 400
rect 23381 368 27000 370
rect 23381 312 23386 368
rect 23442 312 27000 368
rect 23381 310 27000 312
rect 23381 307 23447 310
rect 26200 280 27000 310
<< via3 >>
rect 6316 26148 6380 26212
rect 14412 24516 14476 24580
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 19380 24304 19444 24308
rect 19380 24248 19394 24304
rect 19394 24248 19444 24304
rect 19380 24244 19444 24248
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 8524 23836 8588 23900
rect 15332 23700 15396 23764
rect 21220 23564 21284 23628
rect 6684 23488 6748 23492
rect 6684 23432 6734 23488
rect 6734 23432 6748 23488
rect 6684 23428 6748 23432
rect 14596 23428 14660 23492
rect 17356 23488 17420 23492
rect 17356 23432 17370 23488
rect 17370 23432 17420 23488
rect 17356 23428 17420 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 22692 23156 22756 23220
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 19196 22476 19260 22540
rect 19932 22340 19996 22404
rect 23612 22400 23676 22404
rect 23612 22344 23662 22400
rect 23662 22344 23676 22400
rect 23612 22340 23676 22344
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 21956 22264 22020 22268
rect 21956 22208 22006 22264
rect 22006 22208 22020 22264
rect 21956 22204 22020 22208
rect 18460 21796 18524 21860
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 19380 21388 19444 21452
rect 20668 21388 20732 21452
rect 16436 21252 16500 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 12572 20980 12636 21044
rect 12388 20708 12452 20772
rect 23428 20844 23492 20908
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 6316 20572 6380 20636
rect 19564 20572 19628 20636
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 15148 20028 15212 20092
rect 19380 20088 19444 20092
rect 19380 20032 19430 20088
rect 19430 20032 19444 20088
rect 19380 20028 19444 20032
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 22324 19484 22388 19548
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 21036 19076 21100 19140
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 8524 17988 8588 18052
rect 22508 17988 22572 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 20668 17852 20732 17916
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 15148 17308 15212 17372
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 15332 16764 15396 16828
rect 21588 16628 21652 16692
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 21956 16280 22020 16284
rect 21956 16224 22006 16280
rect 22006 16224 22020 16280
rect 21956 16220 22020 16224
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 22508 15540 22572 15604
rect 16436 15404 16500 15468
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 14412 15132 14476 15196
rect 23428 14996 23492 15060
rect 14596 14860 14660 14924
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 18460 14316 18524 14380
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 6684 13772 6748 13836
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 19196 13500 19260 13564
rect 19380 13364 19444 13428
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 19564 12548 19628 12612
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 21220 12276 21284 12340
rect 22692 12140 22756 12204
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 20668 11868 20732 11932
rect 23612 11868 23676 11932
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 22508 11188 22572 11252
rect 19932 11052 19996 11116
rect 21036 11052 21100 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 17356 10236 17420 10300
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 20668 9556 20732 9620
rect 21588 9616 21652 9620
rect 21588 9560 21602 9616
rect 21602 9560 21652 9616
rect 21588 9556 21652 9560
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 6315 26212 6381 26213
rect 6315 26148 6316 26212
rect 6380 26148 6381 26212
rect 6315 26147 6381 26148
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 6318 20637 6378 26147
rect 14411 24580 14477 24581
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 6683 23492 6749 23493
rect 6683 23428 6684 23492
rect 6748 23428 6749 23492
rect 6683 23427 6749 23428
rect 6315 20636 6381 20637
rect 6315 20572 6316 20636
rect 6380 20572 6381 20636
rect 6315 20571 6381 20572
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 6686 13837 6746 23427
rect 7944 22880 8264 23904
rect 12944 24512 13264 24528
rect 14411 24516 14412 24580
rect 14476 24516 14477 24580
rect 14411 24515 14477 24516
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 8523 23900 8589 23901
rect 8523 23836 8524 23900
rect 8588 23836 8589 23900
rect 8523 23835 8589 23836
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 8526 18053 8586 23835
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12571 21044 12637 21045
rect 12571 20980 12572 21044
rect 12636 20980 12637 21044
rect 12571 20979 12637 20980
rect 12387 20772 12453 20773
rect 12387 20708 12388 20772
rect 12452 20770 12453 20772
rect 12574 20770 12634 20979
rect 12452 20710 12634 20770
rect 12452 20708 12453 20710
rect 12387 20707 12453 20708
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 8523 18052 8589 18053
rect 8523 17988 8524 18052
rect 8588 17988 8589 18052
rect 8523 17987 8589 17988
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 6683 13836 6749 13837
rect 6683 13772 6684 13836
rect 6748 13772 6749 13836
rect 6683 13771 6749 13772
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 14414 15197 14474 24515
rect 17944 23968 18264 24528
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 19379 24308 19445 24309
rect 19379 24244 19380 24308
rect 19444 24244 19445 24308
rect 19379 24243 19445 24244
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 15331 23764 15397 23765
rect 15331 23700 15332 23764
rect 15396 23700 15397 23764
rect 15331 23699 15397 23700
rect 14595 23492 14661 23493
rect 14595 23428 14596 23492
rect 14660 23428 14661 23492
rect 14595 23427 14661 23428
rect 14411 15196 14477 15197
rect 14411 15132 14412 15196
rect 14476 15132 14477 15196
rect 14411 15131 14477 15132
rect 14598 14925 14658 23427
rect 15147 20092 15213 20093
rect 15147 20028 15148 20092
rect 15212 20028 15213 20092
rect 15147 20027 15213 20028
rect 15150 17373 15210 20027
rect 15147 17372 15213 17373
rect 15147 17308 15148 17372
rect 15212 17308 15213 17372
rect 15147 17307 15213 17308
rect 15334 16829 15394 23699
rect 17355 23492 17421 23493
rect 17355 23428 17356 23492
rect 17420 23428 17421 23492
rect 17355 23427 17421 23428
rect 16435 21316 16501 21317
rect 16435 21252 16436 21316
rect 16500 21252 16501 21316
rect 16435 21251 16501 21252
rect 15331 16828 15397 16829
rect 15331 16764 15332 16828
rect 15396 16764 15397 16828
rect 15331 16763 15397 16764
rect 16438 15469 16498 21251
rect 16435 15468 16501 15469
rect 16435 15404 16436 15468
rect 16500 15404 16501 15468
rect 16435 15403 16501 15404
rect 14595 14924 14661 14925
rect 14595 14860 14596 14924
rect 14660 14860 14661 14924
rect 14595 14859 14661 14860
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 17358 10301 17418 23427
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 19195 22540 19261 22541
rect 19195 22476 19196 22540
rect 19260 22476 19261 22540
rect 19195 22475 19261 22476
rect 18459 21860 18525 21861
rect 18459 21796 18460 21860
rect 18524 21796 18525 21860
rect 18459 21795 18525 21796
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 18462 14381 18522 21795
rect 18459 14380 18525 14381
rect 18459 14316 18460 14380
rect 18524 14316 18525 14380
rect 18459 14315 18525 14316
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 19198 13565 19258 22475
rect 19382 21453 19442 24243
rect 21219 23628 21285 23629
rect 21219 23564 21220 23628
rect 21284 23564 21285 23628
rect 21219 23563 21285 23564
rect 19931 22404 19997 22405
rect 19931 22340 19932 22404
rect 19996 22340 19997 22404
rect 19931 22339 19997 22340
rect 19379 21452 19445 21453
rect 19379 21388 19380 21452
rect 19444 21388 19445 21452
rect 19379 21387 19445 21388
rect 19563 20636 19629 20637
rect 19563 20572 19564 20636
rect 19628 20572 19629 20636
rect 19563 20571 19629 20572
rect 19379 20092 19445 20093
rect 19379 20028 19380 20092
rect 19444 20028 19445 20092
rect 19379 20027 19445 20028
rect 19195 13564 19261 13565
rect 19195 13500 19196 13564
rect 19260 13500 19261 13564
rect 19195 13499 19261 13500
rect 19382 13429 19442 20027
rect 19379 13428 19445 13429
rect 19379 13364 19380 13428
rect 19444 13364 19445 13428
rect 19379 13363 19445 13364
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 19566 12613 19626 20571
rect 19563 12612 19629 12613
rect 19563 12548 19564 12612
rect 19628 12548 19629 12612
rect 19563 12547 19629 12548
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 19934 11117 19994 22339
rect 20667 21452 20733 21453
rect 20667 21388 20668 21452
rect 20732 21388 20733 21452
rect 20667 21387 20733 21388
rect 20670 17917 20730 21387
rect 21035 19140 21101 19141
rect 21035 19076 21036 19140
rect 21100 19076 21101 19140
rect 21035 19075 21101 19076
rect 20667 17916 20733 17917
rect 20667 17852 20668 17916
rect 20732 17852 20733 17916
rect 20667 17851 20733 17852
rect 20667 11932 20733 11933
rect 20667 11868 20668 11932
rect 20732 11868 20733 11932
rect 20667 11867 20733 11868
rect 19931 11116 19997 11117
rect 19931 11052 19932 11116
rect 19996 11052 19997 11116
rect 19931 11051 19997 11052
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17355 10300 17421 10301
rect 17355 10236 17356 10300
rect 17420 10236 17421 10300
rect 17355 10235 17421 10236
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 20670 9621 20730 11867
rect 21038 11117 21098 19075
rect 21222 12341 21282 23563
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22691 23220 22757 23221
rect 22691 23156 22692 23220
rect 22756 23156 22757 23220
rect 22691 23155 22757 23156
rect 21955 22268 22021 22269
rect 21955 22204 21956 22268
rect 22020 22204 22021 22268
rect 21955 22203 22021 22204
rect 21587 16692 21653 16693
rect 21587 16628 21588 16692
rect 21652 16628 21653 16692
rect 21587 16627 21653 16628
rect 21219 12340 21285 12341
rect 21219 12276 21220 12340
rect 21284 12276 21285 12340
rect 21219 12275 21285 12276
rect 21035 11116 21101 11117
rect 21035 11052 21036 11116
rect 21100 11052 21101 11116
rect 21035 11051 21101 11052
rect 21590 9621 21650 16627
rect 21958 16285 22018 22203
rect 22323 19548 22389 19549
rect 22323 19484 22324 19548
rect 22388 19484 22389 19548
rect 22323 19483 22389 19484
rect 21955 16284 22021 16285
rect 21955 16220 21956 16284
rect 22020 16220 22021 16284
rect 21955 16219 22021 16220
rect 22326 12450 22386 19483
rect 22507 18052 22573 18053
rect 22507 17988 22508 18052
rect 22572 17988 22573 18052
rect 22507 17987 22573 17988
rect 22510 15605 22570 17987
rect 22507 15604 22573 15605
rect 22507 15540 22508 15604
rect 22572 15540 22573 15604
rect 22507 15539 22573 15540
rect 22326 12390 22570 12450
rect 22510 11253 22570 12390
rect 22694 12205 22754 23155
rect 22944 22336 23264 23360
rect 23611 22404 23677 22405
rect 23611 22340 23612 22404
rect 23676 22340 23677 22404
rect 23611 22339 23677 22340
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 23427 20908 23493 20909
rect 23427 20844 23428 20908
rect 23492 20844 23493 20908
rect 23427 20843 23493 20844
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 23430 15061 23490 20843
rect 23427 15060 23493 15061
rect 23427 14996 23428 15060
rect 23492 14996 23493 15060
rect 23427 14995 23493 14996
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22691 12204 22757 12205
rect 22691 12140 22692 12204
rect 22756 12140 22757 12204
rect 22691 12139 22757 12140
rect 22944 11456 23264 12480
rect 23614 11933 23674 22339
rect 23611 11932 23677 11933
rect 23611 11868 23612 11932
rect 23676 11868 23677 11932
rect 23611 11867 23677 11868
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22507 11252 22573 11253
rect 22507 11188 22508 11252
rect 22572 11188 22573 11252
rect 22507 11187 22573 11188
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 20667 9620 20733 9621
rect 20667 9556 20668 9620
rect 20732 9556 20733 9620
rect 20667 9555 20733 9556
rect 21587 9620 21653 9621
rect 21587 9556 21588 9620
rect 21652 9556 21653 9620
rect 21587 9555 21653 9556
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1676037725
transform 1 0 21896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1676037725
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1676037725
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1676037725
transform 1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1676037725
transform 1 0 24656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1676037725
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1676037725
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1676037725
transform 1 0 15088 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1676037725
transform 1 0 20240 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _098_
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1676037725
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1676037725
transform 1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 15272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 15732 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 8280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 14536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 15272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 5888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _124_
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1676037725
transform 1 0 2116 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 7084 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 5152 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 5244 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 4600 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 17572 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 3956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 18400 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 3312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 7268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 7820 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 9016 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 5152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 6532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 9292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1676037725
transform 1 0 17204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1676037725
transform 1 0 12144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1676037725
transform 1 0 2668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1676037725
transform 1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1676037725
transform 1 0 5520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1676037725
transform 1 0 20608 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1676037725
transform 1 0 23736 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1676037725
transform 1 0 23736 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1676037725
transform 1 0 23552 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1676037725
transform 1 0 9384 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1676037725
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1676037725
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_259
timestamp 1676037725
transform 1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1676037725
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1676037725
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_217
timestamp 1676037725
transform 1 0 21068 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1676037725
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1676037725
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1676037725
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1676037725
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_258
timestamp 1676037725
transform 1 0 24840 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_208
timestamp 1676037725
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1676037725
transform 1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_118
timestamp 1676037725
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp 1676037725
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_216
timestamp 1676037725
transform 1 0 20976 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_223
timestamp 1676037725
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 1676037725
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_180
timestamp 1676037725
transform 1 0 17664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1676037725
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1676037725
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1676037725
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1676037725
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1676037725
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_211
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_240
timestamp 1676037725
transform 1 0 23184 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_246
timestamp 1676037725
transform 1 0 23736 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1676037725
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1676037725
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_179
timestamp 1676037725
transform 1 0 17572 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1676037725
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_191
timestamp 1676037725
transform 1 0 18676 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1676037725
transform 1 0 19044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1676037725
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1676037725
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1676037725
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1676037725
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_216
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_228
timestamp 1676037725
transform 1 0 22080 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_258
timestamp 1676037725
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1676037725
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_197
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_228
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1676037725
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1676037725
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1676037725
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1676037725
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_175
timestamp 1676037725
transform 1 0 17204 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_183
timestamp 1676037725
transform 1 0 17940 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1676037725
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_160
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_206
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1676037725
transform 1 0 20608 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_250
timestamp 1676037725
transform 1 0 24104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_234
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_240
timestamp 1676037725
transform 1 0 23184 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1676037725
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_106
timestamp 1676037725
transform 1 0 10856 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1676037725
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_142
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_148
timestamp 1676037725
transform 1 0 14720 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_231
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_257
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_94
timestamp 1676037725
transform 1 0 9752 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_124
timestamp 1676037725
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_163
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_171
timestamp 1676037725
transform 1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1676037725
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1676037725
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1676037725
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_90
timestamp 1676037725
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1676037725
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_156
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1676037725
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1676037725
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1676037725
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp 1676037725
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_37
timestamp 1676037725
transform 1 0 4508 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_42
timestamp 1676037725
transform 1 0 4968 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_50
timestamp 1676037725
transform 1 0 5704 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 1676037725
transform 1 0 6348 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1676037725
transform 1 0 6900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1676037725
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_100
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1676037725
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1676037725
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_259
timestamp 1676037725
transform 1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_23
timestamp 1676037725
transform 1 0 3220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_42
timestamp 1676037725
transform 1 0 4968 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_75
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_124
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_142
timestamp 1676037725
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_150
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1676037725
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1676037725
transform 1 0 20884 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_248
timestamp 1676037725
transform 1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1676037725
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1676037725
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1676037725
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1676037725
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_46
timestamp 1676037725
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_58
timestamp 1676037725
transform 1 0 6440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_64
timestamp 1676037725
transform 1 0 6992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_169
timestamp 1676037725
transform 1 0 16652 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_231
timestamp 1676037725
transform 1 0 22356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_260
timestamp 1676037725
transform 1 0 25024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1676037725
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_34
timestamp 1676037725
transform 1 0 4232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1676037725
transform 1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_72
timestamp 1676037725
transform 1 0 7728 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_78
timestamp 1676037725
transform 1 0 8280 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1676037725
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_88
timestamp 1676037725
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1676037725
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_247
timestamp 1676037725
transform 1 0 23828 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_251
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_12
timestamp 1676037725
transform 1 0 2208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_20
timestamp 1676037725
transform 1 0 2944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1676037725
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1676037725
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_44
timestamp 1676037725
transform 1 0 5152 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_50
timestamp 1676037725
transform 1 0 5704 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1676037725
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1676037725
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1676037725
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_74
timestamp 1676037725
transform 1 0 7912 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_107
timestamp 1676037725
transform 1 0 10948 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1676037725
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_36
timestamp 1676037725
transform 1 0 4416 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1676037725
transform 1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_44
timestamp 1676037725
transform 1 0 5152 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_50
timestamp 1676037725
transform 1 0 5704 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1676037725
transform 1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_78
timestamp 1676037725
transform 1 0 8280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_83
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1676037725
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1676037725
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1676037725
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1676037725
transform 1 0 7360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 1676037725
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_174
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_216
timestamp 1676037725
transform 1 0 20976 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1676037725
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_34
timestamp 1676037725
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_40
timestamp 1676037725
transform 1 0 4784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_128
timestamp 1676037725
transform 1 0 12880 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_134
timestamp 1676037725
transform 1 0 13432 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1676037725
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_242
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1676037725
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_54
timestamp 1676037725
transform 1 0 6072 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp 1676037725
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_90
timestamp 1676037725
transform 1 0 9384 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1676037725
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_187
timestamp 1676037725
transform 1 0 18308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_202
timestamp 1676037725
transform 1 0 19688 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_229
timestamp 1676037725
transform 1 0 22172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 1676037725
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_17
timestamp 1676037725
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_63
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1676037725
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_128
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_152
timestamp 1676037725
transform 1 0 15088 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1676037725
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_229
timestamp 1676037725
transform 1 0 22172 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_264
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_35
timestamp 1676037725
transform 1 0 4324 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_42
timestamp 1676037725
transform 1 0 4968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_92
timestamp 1676037725
transform 1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1676037725
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_123
timestamp 1676037725
transform 1 0 12420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_131
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1676037725
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1676037725
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_150
timestamp 1676037725
transform 1 0 14904 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_171
timestamp 1676037725
transform 1 0 16836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_175
timestamp 1676037725
transform 1 0 17204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_185
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_208
timestamp 1676037725
transform 1 0 20240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1676037725
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_17
timestamp 1676037725
transform 1 0 2668 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1676037725
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1676037725
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_131
timestamp 1676037725
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1676037725
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1676037725
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_184
timestamp 1676037725
transform 1 0 18032 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1676037725
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_216
timestamp 1676037725
transform 1 0 20976 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_236
timestamp 1676037725
transform 1 0 22816 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_246
timestamp 1676037725
transform 1 0 23736 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1676037725
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1676037725
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1676037725
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_146
timestamp 1676037725
transform 1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_242
timestamp 1676037725
transform 1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1676037725
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_17
timestamp 1676037725
transform 1 0 2668 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1676037725
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_139
timestamp 1676037725
transform 1 0 13892 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1676037725
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_208
timestamp 1676037725
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_248
timestamp 1676037725
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_147
timestamp 1676037725
transform 1 0 14628 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_158
timestamp 1676037725
transform 1 0 15640 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_173
timestamp 1676037725
transform 1 0 17020 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1676037725
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_242
timestamp 1676037725
transform 1 0 23368 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 9384 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 8648 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 17664 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 3956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 17296 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 3312 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1676037725
transform 1 0 10304 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 6072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1676037725
transform 1 0 20792 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 22448 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1676037725
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1676037725
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 7268 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 9844 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 11684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 2760 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16928 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20424 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21528 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20516 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18400 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17848 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13524 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10672 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__159 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__165
timestamp 1676037725
transform 1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21344 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__134
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__139
timestamp 1676037725
transform 1 0 18768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__140
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__162
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__164
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__166
timestamp 1676037725
transform 1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__167
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__132
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__133
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__135
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__136
timestamp 1676037725
transform 1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__137
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__138
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__141
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17296 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__147
timestamp 1676037725
transform 1 0 24104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18952 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__157
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17204 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13984 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__142
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__143
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16008 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__144
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__145
timestamp 1676037725
transform 1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__146
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__148
timestamp 1676037725
transform 1 0 8464 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__149
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__150
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 13064 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13340 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset_top_in
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable_top_in
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal2 6762 1588 6762 1588 0 ccff_head
rlabel metal3 24894 340 24894 340 0 ccff_tail
rlabel metal1 20332 8466 20332 8466 0 chanx_right_in[0]
rlabel metal2 17250 16184 17250 16184 0 chanx_right_in[10]
rlabel metal1 13662 17544 13662 17544 0 chanx_right_in[11]
rlabel metal1 19734 17000 19734 17000 0 chanx_right_in[12]
rlabel metal3 17204 18904 17204 18904 0 chanx_right_in[13]
rlabel metal3 13708 17136 13708 17136 0 chanx_right_in[14]
rlabel metal1 4048 17170 4048 17170 0 chanx_right_in[15]
rlabel metal1 17894 10676 17894 10676 0 chanx_right_in[16]
rlabel metal3 22724 20060 22724 20060 0 chanx_right_in[17]
rlabel metal2 17342 19924 17342 19924 0 chanx_right_in[18]
rlabel metal3 16468 22372 16468 22372 0 chanx_right_in[19]
rlabel metal1 18952 13158 18952 13158 0 chanx_right_in[1]
rlabel metal2 21206 22780 21206 22780 0 chanx_right_in[20]
rlabel metal2 19550 9350 19550 9350 0 chanx_right_in[21]
rlabel metal3 23069 11628 23069 11628 0 chanx_right_in[22]
rlabel metal1 17664 10642 17664 10642 0 chanx_right_in[23]
rlabel metal1 18078 13362 18078 13362 0 chanx_right_in[24]
rlabel metal2 15870 12019 15870 12019 0 chanx_right_in[25]
rlabel metal1 14674 11764 14674 11764 0 chanx_right_in[26]
rlabel metal1 12926 13940 12926 13940 0 chanx_right_in[27]
rlabel metal1 12880 14586 12880 14586 0 chanx_right_in[28]
rlabel metal3 13340 15096 13340 15096 0 chanx_right_in[29]
rlabel metal1 22264 6766 22264 6766 0 chanx_right_in[2]
rlabel metal1 21942 11118 21942 11118 0 chanx_right_in[3]
rlabel metal2 15686 14790 15686 14790 0 chanx_right_in[4]
rlabel metal1 24472 18258 24472 18258 0 chanx_right_in[5]
rlabel metal2 25346 15215 25346 15215 0 chanx_right_in[6]
rlabel metal3 17204 15368 17204 15368 0 chanx_right_in[7]
rlabel metal2 19274 17017 19274 17017 0 chanx_right_in[8]
rlabel via2 19458 16779 19458 16779 0 chanx_right_in[9]
rlabel metal2 25070 1853 25070 1853 0 chanx_right_out[0]
rlabel metal1 24104 5270 24104 5270 0 chanx_right_out[10]
rlabel metal2 24794 4641 24794 4641 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal1 24104 6358 24104 6358 0 chanx_right_out[13]
rlabel metal2 24702 5797 24702 5797 0 chanx_right_out[14]
rlabel metal1 24380 6834 24380 6834 0 chanx_right_out[15]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[16]
rlabel metal3 25584 7684 25584 7684 0 chanx_right_out[17]
rlabel metal1 24426 7922 24426 7922 0 chanx_right_out[18]
rlabel metal1 24104 8534 24104 8534 0 chanx_right_out[19]
rlabel metal3 24250 1156 24250 1156 0 chanx_right_out[1]
rlabel metal2 24702 8109 24702 8109 0 chanx_right_out[20]
rlabel metal1 24426 9010 24426 9010 0 chanx_right_out[21]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[22]
rlabel metal2 24610 9265 24610 9265 0 chanx_right_out[23]
rlabel metal1 24104 10710 24104 10710 0 chanx_right_out[24]
rlabel metal2 24794 10217 24794 10217 0 chanx_right_out[25]
rlabel metal1 24426 11186 24426 11186 0 chanx_right_out[26]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[27]
rlabel metal2 24702 11373 24702 11373 0 chanx_right_out[28]
rlabel metal3 25584 12580 25584 12580 0 chanx_right_out[29]
rlabel metal2 22218 2805 22218 2805 0 chanx_right_out[2]
rlabel metal1 20838 2346 20838 2346 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 25676 3196 25676 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal2 25162 3553 25162 3553 0 chanx_right_out[8]
rlabel metal3 25676 4420 25676 4420 0 chanx_right_out[9]
rlabel metal2 12650 24497 12650 24497 0 chany_top_in[0]
rlabel metal1 16284 19346 16284 19346 0 chany_top_in[10]
rlabel metal2 16974 23324 16974 23324 0 chany_top_in[11]
rlabel metal2 18538 22984 18538 22984 0 chany_top_in[12]
rlabel metal2 17618 24684 17618 24684 0 chany_top_in[13]
rlabel metal1 15778 22542 15778 22542 0 chany_top_in[14]
rlabel metal2 18952 21692 18952 21692 0 chany_top_in[15]
rlabel metal1 16560 21998 16560 21998 0 chany_top_in[16]
rlabel metal2 18998 25493 18998 25493 0 chany_top_in[17]
rlabel metal1 6026 19414 6026 19414 0 chany_top_in[18]
rlabel metal2 16698 18836 16698 18836 0 chany_top_in[19]
rlabel metal1 3956 18734 3956 18734 0 chany_top_in[1]
rlabel metal2 20155 26316 20155 26316 0 chany_top_in[20]
rlabel metal2 20286 26248 20286 26248 0 chany_top_in[21]
rlabel metal4 18492 18088 18492 18088 0 chany_top_in[22]
rlabel metal2 13846 14280 13846 14280 0 chany_top_in[23]
rlabel metal1 5336 18258 5336 18258 0 chany_top_in[24]
rlabel metal4 12604 20876 12604 20876 0 chany_top_in[25]
rlabel metal1 2208 18734 2208 18734 0 chany_top_in[26]
rlabel metal2 21022 22253 21022 22253 0 chany_top_in[27]
rlabel metal2 20102 10659 20102 10659 0 chany_top_in[28]
rlabel metal3 18975 13532 18975 13532 0 chany_top_in[29]
rlabel metal2 6394 19159 6394 19159 0 chany_top_in[2]
rlabel metal1 14214 19822 14214 19822 0 chany_top_in[3]
rlabel metal2 13938 25517 13938 25517 0 chany_top_in[4]
rlabel metal2 14306 25211 14306 25211 0 chany_top_in[5]
rlabel metal2 2070 19686 2070 19686 0 chany_top_in[6]
rlabel metal2 15088 23188 15088 23188 0 chany_top_in[7]
rlabel metal3 18262 21012 18262 21012 0 chany_top_in[8]
rlabel metal2 22034 24174 22034 24174 0 chany_top_in[9]
rlabel metal1 1978 19278 1978 19278 0 chany_top_out[0]
rlabel metal1 4554 23766 4554 23766 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal2 6118 24184 6118 24184 0 chany_top_out[12]
rlabel metal1 4876 24242 4876 24242 0 chany_top_out[13]
rlabel metal1 6946 21012 6946 21012 0 chany_top_out[14]
rlabel metal1 7498 21454 7498 21454 0 chany_top_out[15]
rlabel metal1 6716 23766 6716 23766 0 chany_top_out[16]
rlabel metal1 6578 23188 6578 23188 0 chany_top_out[17]
rlabel metal2 8326 24184 8326 24184 0 chany_top_out[18]
rlabel metal1 7268 24106 7268 24106 0 chany_top_out[19]
rlabel metal2 2070 24218 2070 24218 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8234 23188 8234 23188 0 chany_top_out[21]
rlabel metal1 8970 24242 8970 24242 0 chany_top_out[22]
rlabel metal1 9660 23766 9660 23766 0 chany_top_out[23]
rlabel metal2 10534 24728 10534 24728 0 chany_top_out[24]
rlabel metal2 10902 25034 10902 25034 0 chany_top_out[25]
rlabel metal2 11040 24242 11040 24242 0 chany_top_out[26]
rlabel metal1 11914 23154 11914 23154 0 chany_top_out[27]
rlabel metal2 12282 24973 12282 24973 0 chany_top_out[28]
rlabel metal1 12650 24242 12650 24242 0 chany_top_out[29]
rlabel metal2 2714 23936 2714 23936 0 chany_top_out[2]
rlabel metal1 3220 26418 3220 26418 0 chany_top_out[3]
rlabel metal2 3029 26316 3029 26316 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal1 4324 20978 4324 20978 0 chany_top_out[6]
rlabel metal1 4140 22678 4140 22678 0 chany_top_out[7]
rlabel metal1 3956 23154 3956 23154 0 chany_top_out[8]
rlabel metal1 5060 21454 5060 21454 0 chany_top_out[9]
rlabel metal1 13018 18360 13018 18360 0 clknet_0_prog_clk
rlabel metal1 10534 13158 10534 13158 0 clknet_3_0__leaf_prog_clk
rlabel metal1 17526 12614 17526 12614 0 clknet_3_1__leaf_prog_clk
rlabel metal1 12650 20944 12650 20944 0 clknet_3_2__leaf_prog_clk
rlabel metal2 13570 20162 13570 20162 0 clknet_3_3__leaf_prog_clk
rlabel metal2 16882 15810 16882 15810 0 clknet_3_4__leaf_prog_clk
rlabel via1 21942 13277 21942 13277 0 clknet_3_5__leaf_prog_clk
rlabel metal1 18032 21522 18032 21522 0 clknet_3_6__leaf_prog_clk
rlabel metal1 21804 23290 21804 23290 0 clknet_3_7__leaf_prog_clk
rlabel metal2 6854 5746 6854 5746 0 net1
rlabel metal2 13202 15028 13202 15028 0 net10
rlabel metal1 23920 3026 23920 3026 0 net100
rlabel metal1 22586 4590 22586 4590 0 net101
rlabel metal2 1978 21148 1978 21148 0 net102
rlabel metal2 15962 22831 15962 22831 0 net103
rlabel metal2 17066 23783 17066 23783 0 net104
rlabel metal1 6164 17850 6164 17850 0 net105
rlabel metal1 4048 19482 4048 19482 0 net106
rlabel metal1 7728 17850 7728 17850 0 net107
rlabel metal1 8464 17306 8464 17306 0 net108
rlabel metal1 14812 22134 14812 22134 0 net109
rlabel metal2 14582 23987 14582 23987 0 net11
rlabel metal2 18722 21913 18722 21913 0 net110
rlabel metal2 13754 23885 13754 23885 0 net111
rlabel metal2 15502 24480 15502 24480 0 net112
rlabel metal2 3726 18700 3726 18700 0 net113
rlabel metal1 6348 17306 6348 17306 0 net114
rlabel metal1 7728 18394 7728 18394 0 net115
rlabel metal1 5152 19890 5152 19890 0 net116
rlabel metal1 6946 19482 6946 19482 0 net117
rlabel metal1 4554 18224 4554 18224 0 net118
rlabel metal1 1886 20502 1886 20502 0 net119
rlabel metal1 14398 19754 14398 19754 0 net12
rlabel metal1 9246 20502 9246 20502 0 net120
rlabel metal2 11730 23018 11730 23018 0 net121
rlabel metal1 4324 23086 4324 23086 0 net122
rlabel metal2 12558 24225 12558 24225 0 net123
rlabel metal1 2254 20944 2254 20944 0 net124
rlabel metal1 4462 20434 4462 20434 0 net125
rlabel metal1 2507 21998 2507 21998 0 net126
rlabel metal1 2990 21556 2990 21556 0 net127
rlabel metal1 5796 18122 5796 18122 0 net128
rlabel metal1 4830 18156 4830 18156 0 net129
rlabel metal1 15916 20434 15916 20434 0 net13
rlabel metal2 3634 22610 3634 22610 0 net130
rlabel metal2 13478 21709 13478 21709 0 net131
rlabel metal1 21597 15470 21597 15470 0 net132
rlabel metal1 19366 14382 19366 14382 0 net133
rlabel metal2 20746 24616 20746 24616 0 net134
rlabel metal1 17940 13906 17940 13906 0 net135
rlabel metal1 18630 12682 18630 12682 0 net136
rlabel metal1 21850 11730 21850 11730 0 net137
rlabel metal2 25070 8636 25070 8636 0 net138
rlabel metal1 19136 16218 19136 16218 0 net139
rlabel metal1 15318 20774 15318 20774 0 net14
rlabel metal2 14950 17680 14950 17680 0 net140
rlabel metal2 19826 20366 19826 20366 0 net141
rlabel metal1 14582 20910 14582 20910 0 net142
rlabel metal2 12466 21828 12466 21828 0 net143
rlabel metal1 4968 16966 4968 16966 0 net144
rlabel metal1 10258 20774 10258 20774 0 net145
rlabel metal1 9108 19822 9108 19822 0 net146
rlabel metal1 19918 21624 19918 21624 0 net147
rlabel metal1 9752 19142 9752 19142 0 net148
rlabel metal1 12650 20570 12650 20570 0 net149
rlabel metal1 16284 21862 16284 21862 0 net15
rlabel metal1 11914 18326 11914 18326 0 net150
rlabel metal2 11086 16966 11086 16966 0 net151
rlabel metal1 16744 24378 16744 24378 0 net152
rlabel metal2 10994 16422 10994 16422 0 net153
rlabel metal1 13340 14586 13340 14586 0 net154
rlabel metal2 14122 15538 14122 15538 0 net155
rlabel metal2 16698 17000 16698 17000 0 net156
rlabel metal1 14214 18904 14214 18904 0 net157
rlabel metal1 14352 23698 14352 23698 0 net158
rlabel metal2 20838 20842 20838 20842 0 net159
rlabel metal1 17112 19754 17112 19754 0 net16
rlabel metal2 18906 13583 18906 13583 0 net160
rlabel metal1 21574 22950 21574 22950 0 net161
rlabel metal1 24518 12410 24518 12410 0 net162
rlabel metal2 25070 13600 25070 13600 0 net163
rlabel metal1 22908 7990 22908 7990 0 net164
rlabel metal4 15180 18700 15180 18700 0 net165
rlabel metal1 23966 12750 23966 12750 0 net166
rlabel metal1 21482 16218 21482 16218 0 net167
rlabel metal2 16882 14892 16882 14892 0 net17
rlabel metal1 16468 11322 16468 11322 0 net18
rlabel metal3 17273 13396 17273 13396 0 net19
rlabel metal1 14720 17170 14720 17170 0 net2
rlabel metal3 17043 12580 17043 12580 0 net20
rlabel metal1 19826 22032 19826 22032 0 net21
rlabel metal2 13938 14450 13938 14450 0 net22
rlabel metal1 12006 14552 12006 14552 0 net23
rlabel metal1 22034 6664 22034 6664 0 net24
rlabel metal3 20884 12444 20884 12444 0 net25
rlabel metal1 19826 16048 19826 16048 0 net26
rlabel metal2 17250 17714 17250 17714 0 net27
rlabel metal2 25162 15504 25162 15504 0 net28
rlabel via2 16790 20859 16790 20859 0 net29
rlabel metal3 12650 19652 12650 19652 0 net3
rlabel metal1 18492 17850 18492 17850 0 net30
rlabel metal1 16008 14042 16008 14042 0 net31
rlabel metal1 13386 21420 13386 21420 0 net32
rlabel metal1 16514 19414 16514 19414 0 net33
rlabel metal1 21620 15402 21620 15402 0 net34
rlabel metal2 21758 16150 21758 16150 0 net35
rlabel metal2 16238 17748 16238 17748 0 net36
rlabel metal1 17342 14790 17342 14790 0 net37
rlabel metal1 15134 15130 15134 15130 0 net38
rlabel metal2 20838 18989 20838 18989 0 net39
rlabel metal1 15916 17170 15916 17170 0 net4
rlabel metal2 9062 16439 9062 16439 0 net40
rlabel metal2 6302 17833 6302 17833 0 net41
rlabel metal3 17204 17544 17204 17544 0 net42
rlabel metal1 5543 12274 5543 12274 0 net43
rlabel metal2 4554 16813 4554 16813 0 net44
rlabel metal2 19366 19023 19366 19023 0 net45
rlabel via2 7130 17765 7130 17765 0 net46
rlabel metal1 13340 14042 13340 14042 0 net47
rlabel metal3 17204 20400 17204 20400 0 net48
rlabel metal4 16468 18360 16468 18360 0 net49
rlabel metal2 17342 17527 17342 17527 0 net5
rlabel metal1 2070 18938 2070 18938 0 net50
rlabel metal3 17756 22916 17756 22916 0 net51
rlabel metal1 19504 10234 19504 10234 0 net52
rlabel metal2 18078 9469 18078 9469 0 net53
rlabel metal1 9499 11322 9499 11322 0 net54
rlabel metal1 21574 13906 21574 13906 0 net55
rlabel via2 24518 13821 24518 13821 0 net56
rlabel metal1 19918 15402 19918 15402 0 net57
rlabel via2 20930 18275 20930 18275 0 net58
rlabel metal2 13846 16541 13846 16541 0 net59
rlabel metal2 17894 19465 17894 19465 0 net6
rlabel metal1 18814 18598 18814 18598 0 net60
rlabel metal1 25162 14314 25162 14314 0 net61
rlabel metal1 12013 8874 12013 8874 0 net62
rlabel metal2 18078 19057 18078 19057 0 net63
rlabel metal2 20838 21471 20838 21471 0 net64
rlabel metal1 20884 18394 20884 18394 0 net65
rlabel metal1 20056 19414 20056 19414 0 net66
rlabel metal1 15732 21454 15732 21454 0 net67
rlabel metal1 17894 19754 17894 19754 0 net68
rlabel metal1 18630 18258 18630 18258 0 net69
rlabel metal2 15594 18207 15594 18207 0 net7
rlabel metal1 14628 18598 14628 18598 0 net70
rlabel metal2 23046 9792 23046 9792 0 net71
rlabel metal1 19734 3026 19734 3026 0 net72
rlabel metal2 22218 11084 22218 11084 0 net73
rlabel metal1 23414 4114 23414 4114 0 net74
rlabel metal1 22862 5610 22862 5610 0 net75
rlabel metal1 22310 6358 22310 6358 0 net76
rlabel metal1 22218 5236 22218 5236 0 net77
rlabel metal1 22678 6800 22678 6800 0 net78
rlabel metal1 22770 7378 22770 7378 0 net79
rlabel metal3 13524 17000 13524 17000 0 net8
rlabel metal1 24334 6290 24334 6290 0 net80
rlabel metal1 22862 7820 22862 7820 0 net81
rlabel metal1 22310 8432 22310 8432 0 net82
rlabel metal1 20746 3502 20746 3502 0 net83
rlabel metal1 23690 7378 23690 7378 0 net84
rlabel metal2 22678 8500 22678 8500 0 net85
rlabel metal1 22126 9588 22126 9588 0 net86
rlabel metal1 23184 8466 23184 8466 0 net87
rlabel metal1 22126 10676 22126 10676 0 net88
rlabel metal2 23966 9758 23966 9758 0 net89
rlabel metal2 18630 13804 18630 13804 0 net9
rlabel metal1 22678 11152 22678 11152 0 net90
rlabel metal1 22126 11696 22126 11696 0 net91
rlabel metal2 23966 10982 23966 10982 0 net92
rlabel metal2 23506 10166 23506 10166 0 net93
rlabel metal1 20746 4114 20746 4114 0 net94
rlabel metal2 20930 14144 20930 14144 0 net95
rlabel metal1 22862 2346 22862 2346 0 net96
rlabel metal2 22310 3196 22310 3196 0 net97
rlabel metal1 23782 3502 23782 3502 0 net98
rlabel metal1 22540 4114 22540 4114 0 net99
rlabel metal1 17204 16082 17204 16082 0 prog_clk
rlabel metal2 24518 25238 24518 25238 0 prog_reset_top_in
rlabel metal1 24978 23766 24978 23766 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21390 24242 21390 24242 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 20654 23732 20654 23732 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 22908 22134 22908 22134 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 15134 16626 15134 16626 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal1 18722 19312 18722 19312 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal2 17710 20757 17710 20757 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 25254 19516 25254 19516 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal1 21850 17816 21850 17816 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal1 25300 19482 25300 19482 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal2 20838 17442 20838 17442 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel metal2 22862 19380 22862 19380 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 23966 15470 23966 15470 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 22908 17714 22908 17714 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal1 23322 12274 23322 12274 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24886 15130 24886 15130 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal1 23000 12954 23000 12954 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal1 24058 12376 24058 12376 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal2 21022 21624 21022 21624 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 20700 20978 20700 20978 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 21298 13804 21298 13804 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 20194 13362 20194 13362 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 21114 16762 21114 16762 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 20233 16762 20233 16762 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal1 20102 16422 20102 16422 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal2 20194 17952 20194 17952 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal2 18630 14620 18630 14620 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal2 18814 17306 18814 17306 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal1 23131 21318 23131 21318 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal2 17526 23868 17526 23868 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17710 13804 17710 13804 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18308 14518 18308 14518 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 20838 12716 20838 12716 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 19826 17714 19826 17714 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20424 12070 20424 12070 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal1 20417 12410 20417 12410 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal1 20240 15538 20240 15538 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 23092 20978 23092 20978 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal2 21850 23766 21850 23766 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal2 16422 24412 16422 24412 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal1 15916 18666 15916 18666 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal2 14950 19550 14950 19550 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 14950 22746 14950 22746 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel metal1 15226 20230 15226 20230 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal2 15042 21114 15042 21114 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 12650 21488 12650 21488 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal1 14536 19482 14536 19482 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 12282 22066 12282 22066 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal1 13294 21114 13294 21114 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 10672 20978 10672 20978 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal1 14030 22066 14030 22066 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 9614 19890 9614 19890 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel via2 14398 19907 14398 19907 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 18538 21012 18538 21012 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal1 17756 20366 17756 20366 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 11040 17306 11040 17306 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal1 13386 18632 13386 18632 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 13478 18156 13478 18156 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel metal1 15364 19414 15364 19414 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 12926 16422 12926 16422 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal1 14352 17782 14352 17782 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 12006 14892 12006 14892 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal1 14858 16218 14858 16218 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 18676 23630 18676 23630 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal1 20746 22508 20746 22508 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 11270 15572 11270 15572 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal1 13340 14926 13340 14926 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 14168 13226 14168 13226 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 15502 13498 15502 13498 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14582 14178 14582 14178 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal1 17526 13430 17526 13430 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16284 14518 16284 14518 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 16284 23630 16284 23630 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal2 19550 23018 19550 23018 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 15410 22950 15410 22950 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 21758 9758 21758 9758 0 sb_0__0_.mux_right_track_0.out
rlabel metal1 19550 21352 19550 21352 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22402 19856 22402 19856 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22034 19448 22034 19448 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 24610 11424 24610 11424 0 sb_0__0_.mux_right_track_10.out
rlabel metal2 24610 19754 24610 19754 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24610 11118 24610 11118 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24518 8058 24518 8058 0 sb_0__0_.mux_right_track_12.out
rlabel via3 22011 16252 22011 16252 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 7854 24104 7854 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20792 9350 20792 9350 0 sb_0__0_.mux_right_track_14.out
rlabel metal1 24150 16218 24150 16218 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21758 9520 21758 9520 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20194 7854 20194 7854 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 24150 14314 24150 14314 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19872 12852 19872 12852 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20194 9996 20194 9996 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 24978 13362 24978 13362 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20424 10642 20424 10642 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19136 9078 19136 9078 0 sb_0__0_.mux_right_track_2.out
rlabel metal1 24610 22406 24610 22406 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23897 9078 23897 9078 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21482 6766 21482 6766 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 21114 13974 21114 13974 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20976 12614 20976 12614 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19090 9010 19090 9010 0 sb_0__0_.mux_right_track_30.out
rlabel metal1 20838 16150 20838 16150 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18952 9554 18952 9554 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 8840 24702 8840 0 sb_0__0_.mux_right_track_32.out
rlabel metal1 21206 15572 21206 15572 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22402 8942 22402 8942 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24518 5678 24518 5678 0 sb_0__0_.mux_right_track_34.out
rlabel metal1 19734 14246 19734 14246 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20332 14518 20332 14518 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 21735 16660 21735 16660 0 sb_0__0_.mux_right_track_4.out
rlabel metal2 25070 23936 25070 23936 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22034 17136 22034 17136 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24518 6766 24518 6766 0 sb_0__0_.mux_right_track_44.out
rlabel metal1 17618 14042 17618 14042 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 14042 17158 14042 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24472 4590 24472 4590 0 sb_0__0_.mux_right_track_46.out
rlabel metal1 20332 12954 20332 12954 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20470 8534 20470 8534 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23828 3570 23828 3570 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 21390 12138 21390 12138 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21482 9724 21482 9724 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 2414 24058 2414 0 sb_0__0_.mux_right_track_50.out
rlabel metal1 25116 9894 25116 9894 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23414 10098 23414 10098 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12742 10642 12742 10642 0 sb_0__0_.mux_right_track_6.out
rlabel metal2 19458 23341 19458 23341 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24978 19499 24978 19499 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10304 15470 10304 15470 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21114 10166 21114 10166 0 sb_0__0_.mux_right_track_8.out
rlabel metal1 20700 18190 20700 18190 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 10030 24104 10030 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 12558 16507 12558 16507 0 sb_0__0_.mux_top_track_0.out
rlabel metal1 14858 18938 14858 18938 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15686 19482 15686 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 19482 14904 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9108 21862 9108 21862 0 sb_0__0_.mux_top_track_10.out
rlabel metal1 14766 21012 14766 21012 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14306 21301 14306 21301 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 4738 20604 4738 20604 0 sb_0__0_.mux_top_track_12.out
rlabel metal1 15042 19958 15042 19958 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4922 21964 4922 21964 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8188 17782 8188 17782 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 15824 21862 15824 21862 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10626 22746 10626 22746 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6854 20230 6854 20230 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 14720 21114 14720 21114 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 6026 20655 6026 20655 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6118 18428 6118 18428 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 10396 19822 10396 19822 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6026 19788 6026 19788 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6486 23086 6486 23086 0 sb_0__0_.mux_top_track_2.out
rlabel metal1 19458 21930 19458 21930 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15594 22066 15594 22066 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8188 17170 8188 17170 0 sb_0__0_.mux_top_track_28.out
rlabel metal2 12098 18870 12098 18870 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7406 19380 7406 19380 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7866 17646 7866 17646 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 16376 20026 16376 20026 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7958 19380 7958 19380 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4370 19380 4370 19380 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 14720 18122 14720 18122 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11224 18054 11224 18054 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6394 17646 6394 17646 0 sb_0__0_.mux_top_track_34.out
rlabel metal1 15594 17068 15594 17068 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9936 16966 9936 16966 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9890 22202 9890 22202 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 20102 22746 20102 22746 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10166 22610 10166 22610 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5014 19108 5014 19108 0 sb_0__0_.mux_top_track_44.out
rlabel via2 15594 15963 15594 15963 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7406 19822 7406 19822 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6624 18258 6624 18258 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 14904 15334 14904 15334 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12098 15810 12098 15810 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7590 19142 7590 19142 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 19458 16184 19458 16184 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13938 15776 13938 15776 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5796 18734 5796 18734 0 sb_0__0_.mux_top_track_50.out
rlabel metal1 15456 17306 15456 17306 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13386 18054 13386 18054 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6854 24038 6854 24038 0 sb_0__0_.mux_top_track_6.out
rlabel metal1 15778 21658 15778 21658 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18952 22746 18952 22746 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15594 23528 15594 23528 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 1610 20332 1610 20332 0 sb_0__0_.mux_top_track_8.out
rlabel metal1 17204 22746 17204 22746 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4186 24004 4186 24004 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 820 22644 820 22644 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 820 23732 820 23732 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 3772 21998 3772 21998 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 2231 21590 2231 21590 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
