magic
tech sky130A
magscale 1 2
timestamp 1682556457
<< viali >>
rect 18981 54281 19015 54315
rect 18153 54213 18187 54247
rect 2237 54145 2271 54179
rect 4169 54145 4203 54179
rect 6745 54145 6779 54179
rect 13737 54145 13771 54179
rect 14105 54145 14139 54179
rect 15117 54145 15151 54179
rect 15393 54145 15427 54179
rect 17049 54145 17083 54179
rect 17325 54145 17359 54179
rect 17877 54145 17911 54179
rect 19717 54145 19751 54179
rect 21189 54145 21223 54179
rect 22293 54145 22327 54179
rect 23397 54145 23431 54179
rect 24593 54145 24627 54179
rect 2513 54077 2547 54111
rect 4445 54077 4479 54111
rect 7113 54077 7147 54111
rect 19441 54077 19475 54111
rect 21373 54009 21407 54043
rect 21925 54009 21959 54043
rect 25237 54009 25271 54043
rect 13553 53941 13587 53975
rect 14933 53941 14967 53975
rect 16865 53941 16899 53975
rect 17693 53941 17727 53975
rect 22937 53941 22971 53975
rect 24041 53941 24075 53975
rect 25237 53737 25271 53771
rect 24225 53669 24259 53703
rect 2053 53601 2087 53635
rect 5733 53601 5767 53635
rect 1777 53533 1811 53567
rect 5457 53533 5491 53567
rect 22109 53533 22143 53567
rect 22385 53533 22419 53567
rect 23121 53533 23155 53567
rect 24593 53533 24627 53567
rect 22569 53397 22603 53431
rect 23765 53397 23799 53431
rect 4997 53193 5031 53227
rect 6561 53193 6595 53227
rect 25237 53193 25271 53227
rect 22477 53125 22511 53159
rect 22845 53125 22879 53159
rect 5181 53057 5215 53091
rect 6745 53057 6779 53091
rect 23489 53057 23523 53091
rect 24593 53057 24627 53091
rect 23029 52921 23063 52955
rect 24133 52853 24167 52887
rect 7665 52649 7699 52683
rect 23121 52649 23155 52683
rect 25329 52649 25363 52683
rect 7849 52445 7883 52479
rect 23305 52445 23339 52479
rect 23765 52445 23799 52479
rect 24685 52445 24719 52479
rect 23949 52309 23983 52343
rect 8861 52105 8895 52139
rect 24961 52037 24995 52071
rect 8769 51969 8803 52003
rect 22937 51969 22971 52003
rect 24133 51969 24167 52003
rect 25237 51901 25271 51935
rect 24317 51833 24351 51867
rect 23581 51765 23615 51799
rect 24133 51561 24167 51595
rect 24593 51561 24627 51595
rect 23857 51493 23891 51527
rect 24041 51289 24075 51323
rect 24961 51289 24995 51323
rect 25053 51221 25087 51255
rect 7941 51017 7975 51051
rect 7481 50881 7515 50915
rect 24593 50881 24627 50915
rect 24961 50881 24995 50915
rect 7573 50677 7607 50711
rect 8401 50677 8435 50711
rect 25053 50677 25087 50711
rect 25513 50133 25547 50167
rect 24501 49793 24535 49827
rect 24777 49725 24811 49759
rect 22569 49181 22603 49215
rect 24777 49113 24811 49147
rect 25145 49113 25179 49147
rect 23213 49045 23247 49079
rect 25237 49045 25271 49079
rect 10517 48841 10551 48875
rect 7941 48773 7975 48807
rect 10977 48773 11011 48807
rect 10057 48705 10091 48739
rect 7757 48637 7791 48671
rect 8401 48637 8435 48671
rect 10149 48501 10183 48535
rect 25421 48501 25455 48535
rect 8309 48229 8343 48263
rect 6561 48161 6595 48195
rect 9137 48093 9171 48127
rect 10276 48093 10310 48127
rect 11472 48093 11506 48127
rect 25145 48093 25179 48127
rect 6837 48025 6871 48059
rect 9781 48025 9815 48059
rect 8585 47957 8619 47991
rect 10379 47957 10413 47991
rect 11575 47957 11609 47991
rect 25237 47957 25271 47991
rect 8861 47685 8895 47719
rect 12484 47617 12518 47651
rect 24869 47617 24903 47651
rect 25329 47617 25363 47651
rect 8677 47549 8711 47583
rect 9321 47549 9355 47583
rect 8401 47413 8435 47447
rect 12587 47413 12621 47447
rect 25145 47413 25179 47447
rect 9781 47209 9815 47243
rect 10333 47209 10367 47243
rect 11069 47209 11103 47243
rect 10701 47141 10735 47175
rect 14289 47073 14323 47107
rect 9137 47005 9171 47039
rect 10241 47005 10275 47039
rect 13312 47005 13346 47039
rect 22661 47005 22695 47039
rect 13415 46937 13449 46971
rect 14473 46937 14507 46971
rect 16129 46937 16163 46971
rect 23305 46937 23339 46971
rect 25421 46869 25455 46903
rect 12357 46597 12391 46631
rect 14657 46597 14691 46631
rect 25329 46529 25363 46563
rect 12173 46461 12207 46495
rect 14013 46461 14047 46495
rect 14473 46461 14507 46495
rect 16313 46461 16347 46495
rect 25145 46325 25179 46359
rect 9781 46121 9815 46155
rect 10793 45985 10827 46019
rect 12081 45985 12115 46019
rect 15761 45985 15795 46019
rect 9137 45917 9171 45951
rect 10609 45917 10643 45951
rect 15577 45917 15611 45951
rect 24869 45917 24903 45951
rect 25329 45917 25363 45951
rect 17417 45849 17451 45883
rect 25145 45781 25179 45815
rect 12173 45577 12207 45611
rect 9505 45509 9539 45543
rect 11713 45441 11747 45475
rect 12541 45441 12575 45475
rect 9321 45373 9355 45407
rect 10977 45373 11011 45407
rect 11805 45237 11839 45271
rect 25421 45237 25455 45271
rect 10885 45033 10919 45067
rect 9137 44897 9171 44931
rect 11345 44829 11379 44863
rect 25329 44829 25363 44863
rect 9413 44761 9447 44795
rect 11989 44761 12023 44795
rect 25145 44693 25179 44727
rect 10885 44489 10919 44523
rect 10241 44353 10275 44387
rect 24777 44353 24811 44387
rect 25145 44353 25179 44387
rect 11253 44285 11287 44319
rect 25329 44217 25363 44251
rect 11621 44149 11655 44183
rect 10609 43945 10643 43979
rect 20821 43809 20855 43843
rect 22569 43809 22603 43843
rect 9965 43741 9999 43775
rect 20545 43741 20579 43775
rect 22293 43605 22327 43639
rect 25513 43605 25547 43639
rect 25145 43333 25179 43367
rect 25237 43061 25271 43095
rect 9952 42857 9986 42891
rect 9689 42721 9723 42755
rect 11989 42721 12023 42755
rect 24777 42585 24811 42619
rect 25145 42585 25179 42619
rect 11437 42517 11471 42551
rect 11713 42517 11747 42551
rect 25237 42517 25271 42551
rect 25421 41973 25455 42007
rect 24777 41497 24811 41531
rect 25145 41497 25179 41531
rect 25237 41429 25271 41463
rect 19441 41089 19475 41123
rect 24225 41089 24259 41123
rect 24685 41089 24719 41123
rect 25329 41089 25363 41123
rect 20085 40885 20119 40919
rect 24501 40885 24535 40919
rect 25145 40885 25179 40919
rect 25329 40477 25363 40511
rect 24685 40341 24719 40375
rect 24869 40341 24903 40375
rect 25145 40341 25179 40375
rect 25145 40069 25179 40103
rect 24593 40001 24627 40035
rect 25329 39865 25363 39899
rect 24409 39797 24443 39831
rect 11897 39593 11931 39627
rect 24777 39593 24811 39627
rect 11253 39389 11287 39423
rect 24225 39321 24259 39355
rect 25145 39321 25179 39355
rect 25329 39321 25363 39355
rect 24501 39253 24535 39287
rect 8585 39049 8619 39083
rect 8769 38913 8803 38947
rect 24225 38913 24259 38947
rect 24685 38913 24719 38947
rect 24041 38709 24075 38743
rect 25329 38709 25363 38743
rect 23857 38437 23891 38471
rect 18245 38301 18279 38335
rect 24041 38301 24075 38335
rect 24593 38301 24627 38335
rect 18889 38165 18923 38199
rect 23489 38165 23523 38199
rect 25237 38165 25271 38199
rect 12357 37961 12391 37995
rect 11713 37825 11747 37859
rect 23029 37825 23063 37859
rect 24041 37825 24075 37859
rect 22753 37757 22787 37791
rect 24961 37689 24995 37723
rect 24685 37621 24719 37655
rect 22293 37213 22327 37247
rect 23397 37213 23431 37247
rect 24593 37213 24627 37247
rect 24041 37145 24075 37179
rect 22937 37077 22971 37111
rect 25237 37077 25271 37111
rect 20545 36873 20579 36907
rect 24225 36873 24259 36907
rect 22293 36737 22327 36771
rect 23581 36737 23615 36771
rect 24685 36737 24719 36771
rect 22937 36533 22971 36567
rect 25329 36533 25363 36567
rect 23949 36329 23983 36363
rect 25237 36329 25271 36363
rect 19993 36125 20027 36159
rect 20637 36125 20671 36159
rect 21097 36125 21131 36159
rect 22201 36125 22235 36159
rect 23305 36125 23339 36159
rect 24593 36125 24627 36159
rect 21741 36057 21775 36091
rect 22845 35989 22879 36023
rect 8769 35785 8803 35819
rect 21097 35785 21131 35819
rect 22477 35785 22511 35819
rect 11713 35717 11747 35751
rect 21189 35717 21223 35751
rect 8953 35649 8987 35683
rect 9413 35649 9447 35683
rect 19625 35649 19659 35683
rect 22385 35649 22419 35683
rect 23213 35649 23247 35683
rect 24317 35649 24351 35683
rect 9689 35581 9723 35615
rect 11161 35581 11195 35615
rect 21281 35581 21315 35615
rect 22569 35581 22603 35615
rect 23857 35513 23891 35547
rect 11621 35445 11655 35479
rect 20269 35445 20303 35479
rect 20729 35445 20763 35479
rect 22017 35445 22051 35479
rect 24961 35445 24995 35479
rect 18705 35241 18739 35275
rect 21741 35173 21775 35207
rect 22109 35173 22143 35207
rect 19349 35105 19383 35139
rect 23213 35105 23247 35139
rect 23305 35105 23339 35139
rect 18889 35037 18923 35071
rect 19625 35037 19659 35071
rect 20729 35037 20763 35071
rect 22293 35037 22327 35071
rect 24593 35037 24627 35071
rect 23121 34969 23155 35003
rect 23949 34969 23983 35003
rect 18245 34901 18279 34935
rect 20269 34901 20303 34935
rect 21373 34901 21407 34935
rect 22753 34901 22787 34935
rect 23765 34901 23799 34935
rect 24133 34901 24167 34935
rect 25237 34901 25271 34935
rect 19165 34697 19199 34731
rect 21373 34697 21407 34731
rect 18061 34561 18095 34595
rect 18521 34561 18555 34595
rect 19625 34561 19659 34595
rect 20269 34561 20303 34595
rect 20729 34561 20763 34595
rect 22017 34561 22051 34595
rect 23121 34561 23155 34595
rect 24225 34561 24259 34595
rect 22661 34493 22695 34527
rect 23765 34493 23799 34527
rect 17877 34357 17911 34391
rect 24869 34357 24903 34391
rect 10425 34153 10459 34187
rect 19704 34153 19738 34187
rect 25237 34153 25271 34187
rect 21189 34085 21223 34119
rect 23397 34085 23431 34119
rect 15117 34017 15151 34051
rect 19441 34017 19475 34051
rect 21649 34017 21683 34051
rect 9781 33949 9815 33983
rect 17049 33949 17083 33983
rect 18153 33949 18187 33983
rect 24041 33949 24075 33983
rect 24593 33949 24627 33983
rect 14381 33881 14415 33915
rect 15577 33881 15611 33915
rect 17693 33881 17727 33915
rect 21925 33881 21959 33915
rect 18797 33813 18831 33847
rect 23857 33813 23891 33847
rect 16221 33609 16255 33643
rect 16497 33609 16531 33643
rect 18153 33609 18187 33643
rect 21281 33609 21315 33643
rect 24685 33609 24719 33643
rect 25329 33609 25363 33643
rect 17509 33473 17543 33507
rect 18613 33473 18647 33507
rect 19073 33473 19107 33507
rect 22017 33473 22051 33507
rect 24593 33473 24627 33507
rect 25421 33473 25455 33507
rect 19533 33405 19567 33439
rect 19809 33405 19843 33439
rect 22293 33405 22327 33439
rect 24777 33405 24811 33439
rect 18889 33269 18923 33303
rect 21649 33269 21683 33303
rect 23765 33269 23799 33303
rect 24225 33269 24259 33303
rect 9321 33065 9355 33099
rect 18429 33065 18463 33099
rect 18705 33065 18739 33099
rect 18981 33065 19015 33099
rect 22556 33065 22590 33099
rect 24041 33065 24075 33099
rect 21189 32997 21223 33031
rect 16037 32929 16071 32963
rect 17233 32929 17267 32963
rect 19717 32929 19751 32963
rect 22293 32929 22327 32963
rect 25053 32929 25087 32963
rect 25145 32929 25179 32963
rect 9505 32861 9539 32895
rect 15761 32861 15795 32895
rect 16957 32861 16991 32895
rect 17785 32861 17819 32895
rect 19441 32861 19475 32895
rect 21833 32861 21867 32895
rect 24961 32861 24995 32895
rect 15853 32793 15887 32827
rect 17049 32793 17083 32827
rect 15393 32725 15427 32759
rect 16589 32725 16623 32759
rect 21649 32725 21683 32759
rect 24593 32725 24627 32759
rect 9045 32521 9079 32555
rect 21281 32521 21315 32555
rect 15393 32453 15427 32487
rect 16865 32453 16899 32487
rect 19901 32453 19935 32487
rect 22017 32453 22051 32487
rect 22753 32453 22787 32487
rect 9229 32385 9263 32419
rect 23397 32385 23431 32419
rect 16129 32317 16163 32351
rect 17693 32317 17727 32351
rect 17969 32317 18003 32351
rect 20637 32317 20671 32351
rect 23673 32317 23707 32351
rect 16681 32181 16715 32215
rect 19441 32181 19475 32215
rect 25145 32181 25179 32215
rect 9873 31977 9907 32011
rect 16037 31977 16071 32011
rect 16681 31977 16715 32011
rect 21189 31977 21223 32011
rect 21465 31977 21499 32011
rect 13553 31909 13587 31943
rect 16497 31909 16531 31943
rect 18797 31909 18831 31943
rect 23857 31909 23891 31943
rect 25237 31909 25271 31943
rect 12357 31841 12391 31875
rect 14289 31841 14323 31875
rect 14565 31841 14599 31875
rect 17049 31841 17083 31875
rect 17325 31841 17359 31875
rect 22569 31841 22603 31875
rect 9229 31773 9263 31807
rect 11713 31773 11747 31807
rect 12909 31773 12943 31807
rect 19441 31773 19475 31807
rect 21649 31773 21683 31807
rect 22477 31773 22511 31807
rect 23213 31773 23247 31807
rect 24593 31773 24627 31807
rect 19717 31705 19751 31739
rect 22017 31637 22051 31671
rect 22385 31637 22419 31671
rect 20637 31433 20671 31467
rect 21557 31433 21591 31467
rect 22661 31433 22695 31467
rect 25145 31433 25179 31467
rect 14013 31365 14047 31399
rect 17049 31365 17083 31399
rect 10517 31297 10551 31331
rect 12265 31297 12299 31331
rect 13369 31297 13403 31331
rect 14565 31297 14599 31331
rect 15669 31297 15703 31331
rect 17325 31297 17359 31331
rect 17969 31297 18003 31331
rect 18429 31297 18463 31331
rect 20729 31297 20763 31331
rect 22017 31297 22051 31331
rect 23397 31297 23431 31331
rect 19625 31229 19659 31263
rect 20821 31229 20855 31263
rect 23673 31229 23707 31263
rect 12909 31161 12943 31195
rect 16313 31161 16347 31195
rect 11161 31093 11195 31127
rect 15209 31093 15243 31127
rect 16773 31093 16807 31127
rect 19073 31093 19107 31127
rect 20269 31093 20303 31127
rect 11253 30889 11287 30923
rect 20361 30889 20395 30923
rect 22845 30889 22879 30923
rect 25237 30889 25271 30923
rect 15945 30821 15979 30855
rect 20085 30821 20119 30855
rect 16497 30753 16531 30787
rect 17141 30753 17175 30787
rect 17417 30753 17451 30787
rect 18889 30753 18923 30787
rect 21097 30753 21131 30787
rect 21373 30753 21407 30787
rect 10609 30685 10643 30719
rect 11713 30685 11747 30719
rect 12817 30685 12851 30719
rect 16405 30685 16439 30719
rect 19441 30685 19475 30719
rect 23305 30685 23339 30719
rect 24593 30685 24627 30719
rect 14289 30617 14323 30651
rect 15025 30617 15059 30651
rect 16313 30617 16347 30651
rect 12357 30549 12391 30583
rect 13461 30549 13495 30583
rect 13829 30549 13863 30583
rect 15577 30549 15611 30583
rect 20545 30549 20579 30583
rect 23949 30549 23983 30583
rect 14381 30345 14415 30379
rect 17325 30345 17359 30379
rect 9689 30277 9723 30311
rect 11161 30277 11195 30311
rect 12909 30277 12943 30311
rect 18705 30277 18739 30311
rect 20361 30277 20395 30311
rect 9045 30209 9079 30243
rect 10517 30209 10551 30243
rect 14841 30209 14875 30243
rect 16405 30209 16439 30243
rect 17233 30209 17267 30243
rect 18061 30209 18095 30243
rect 20269 30209 20303 30243
rect 21189 30209 21223 30243
rect 22109 30209 22143 30243
rect 12633 30141 12667 30175
rect 15577 30141 15611 30175
rect 17417 30141 17451 30175
rect 19165 30141 19199 30175
rect 20453 30141 20487 30175
rect 22753 30141 22787 30175
rect 23029 30141 23063 30175
rect 24961 30141 24995 30175
rect 16313 30073 16347 30107
rect 21373 30073 21407 30107
rect 22293 30073 22327 30107
rect 16037 30005 16071 30039
rect 16865 30005 16899 30039
rect 19901 30005 19935 30039
rect 24501 30005 24535 30039
rect 23949 29733 23983 29767
rect 15577 29665 15611 29699
rect 16497 29665 16531 29699
rect 20085 29665 20119 29699
rect 21097 29665 21131 29699
rect 21189 29665 21223 29699
rect 10149 29597 10183 29631
rect 11253 29597 11287 29631
rect 13737 29597 13771 29631
rect 14565 29597 14599 29631
rect 15393 29597 15427 29631
rect 17141 29597 17175 29631
rect 19809 29597 19843 29631
rect 19901 29597 19935 29631
rect 21005 29597 21039 29631
rect 21925 29597 21959 29631
rect 23305 29597 23339 29631
rect 24593 29597 24627 29631
rect 11529 29529 11563 29563
rect 16129 29529 16163 29563
rect 17417 29529 17451 29563
rect 22661 29529 22695 29563
rect 10793 29461 10827 29495
rect 13001 29461 13035 29495
rect 13553 29461 13587 29495
rect 14381 29461 14415 29495
rect 15025 29461 15059 29495
rect 15485 29461 15519 29495
rect 18889 29461 18923 29495
rect 19441 29461 19475 29495
rect 20637 29461 20671 29495
rect 25237 29461 25271 29495
rect 12633 29257 12667 29291
rect 15117 29257 15151 29291
rect 19993 29257 20027 29291
rect 20085 29257 20119 29291
rect 22477 29257 22511 29291
rect 23673 29257 23707 29291
rect 9689 29189 9723 29223
rect 11713 29189 11747 29223
rect 15853 29189 15887 29223
rect 21465 29189 21499 29223
rect 22385 29189 22419 29223
rect 11989 29121 12023 29155
rect 13093 29121 13127 29155
rect 16865 29121 16899 29155
rect 17957 29121 17991 29155
rect 20821 29121 20855 29155
rect 23581 29121 23615 29155
rect 24409 29121 24443 29155
rect 9413 29053 9447 29087
rect 14841 29053 14875 29087
rect 15945 29053 15979 29087
rect 16129 29053 16163 29087
rect 19349 29053 19383 29087
rect 20269 29053 20303 29087
rect 22661 29053 22695 29087
rect 23765 29053 23799 29087
rect 11161 28985 11195 29019
rect 18613 28985 18647 29019
rect 19625 28985 19659 29019
rect 22017 28985 22051 29019
rect 23213 28985 23247 29019
rect 25053 28985 25087 29019
rect 13356 28917 13390 28951
rect 15485 28917 15519 28951
rect 17509 28917 17543 28951
rect 18889 28917 18923 28951
rect 19165 28917 19199 28951
rect 9689 28713 9723 28747
rect 12817 28713 12851 28747
rect 23857 28713 23891 28747
rect 24133 28713 24167 28747
rect 15485 28645 15519 28679
rect 17877 28645 17911 28679
rect 10241 28577 10275 28611
rect 13553 28577 13587 28611
rect 14749 28577 14783 28611
rect 14841 28577 14875 28611
rect 15945 28577 15979 28611
rect 16037 28577 16071 28611
rect 17233 28577 17267 28611
rect 18521 28577 18555 28611
rect 22753 28577 22787 28611
rect 25053 28577 25087 28611
rect 25145 28577 25179 28611
rect 7941 28509 7975 28543
rect 11069 28509 11103 28543
rect 15853 28509 15887 28543
rect 17049 28509 17083 28543
rect 18337 28509 18371 28543
rect 20821 28509 20855 28543
rect 22661 28509 22695 28543
rect 8585 28441 8619 28475
rect 11345 28441 11379 28475
rect 18245 28441 18279 28475
rect 19441 28441 19475 28475
rect 20177 28441 20211 28475
rect 21557 28441 21591 28475
rect 23213 28441 23247 28475
rect 23397 28441 23431 28475
rect 23673 28441 23707 28475
rect 10057 28373 10091 28407
rect 10149 28373 10183 28407
rect 13185 28373 13219 28407
rect 14289 28373 14323 28407
rect 14657 28373 14691 28407
rect 16681 28373 16715 28407
rect 17141 28373 17175 28407
rect 18889 28373 18923 28407
rect 22201 28373 22235 28407
rect 22569 28373 22603 28407
rect 24593 28373 24627 28407
rect 24961 28373 24995 28407
rect 10425 28169 10459 28203
rect 10701 28169 10735 28203
rect 11253 28169 11287 28203
rect 13553 28169 13587 28203
rect 15761 28169 15795 28203
rect 16957 28169 16991 28203
rect 19349 28169 19383 28203
rect 20453 28169 20487 28203
rect 24961 28169 24995 28203
rect 8677 28033 8711 28067
rect 11805 28033 11839 28067
rect 14013 28033 14047 28067
rect 17601 28033 17635 28067
rect 19809 28033 19843 28067
rect 21005 28033 21039 28067
rect 22017 28033 22051 28067
rect 25053 28033 25087 28067
rect 8953 27965 8987 27999
rect 12081 27965 12115 27999
rect 14289 27965 14323 27999
rect 17877 27965 17911 27999
rect 21189 27965 21223 27999
rect 22293 27965 22327 27999
rect 25145 27965 25179 27999
rect 24593 27897 24627 27931
rect 16129 27829 16163 27863
rect 16405 27829 16439 27863
rect 23765 27829 23799 27863
rect 24133 27829 24167 27863
rect 10136 27625 10170 27659
rect 11897 27625 11931 27659
rect 14565 27625 14599 27659
rect 18613 27625 18647 27659
rect 20900 27625 20934 27659
rect 13737 27557 13771 27591
rect 14197 27557 14231 27591
rect 20085 27557 20119 27591
rect 9873 27489 9907 27523
rect 15485 27489 15519 27523
rect 16589 27489 16623 27523
rect 17785 27489 17819 27523
rect 23397 27489 23431 27523
rect 25145 27489 25179 27523
rect 12633 27421 12667 27455
rect 13093 27421 13127 27455
rect 15209 27421 15243 27455
rect 17601 27421 17635 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 20637 27421 20671 27455
rect 23213 27421 23247 27455
rect 23305 27421 23339 27455
rect 12173 27353 12207 27387
rect 25053 27353 25087 27387
rect 9137 27285 9171 27319
rect 11621 27285 11655 27319
rect 12449 27285 12483 27319
rect 14381 27285 14415 27319
rect 14841 27285 14875 27319
rect 15301 27285 15335 27319
rect 16037 27285 16071 27319
rect 16405 27285 16439 27319
rect 16497 27285 16531 27319
rect 17233 27285 17267 27319
rect 17693 27285 17727 27319
rect 22385 27285 22419 27319
rect 22845 27285 22879 27319
rect 24133 27285 24167 27319
rect 24593 27285 24627 27319
rect 24961 27285 24995 27319
rect 11161 27081 11195 27115
rect 12541 27081 12575 27115
rect 13001 27081 13035 27115
rect 20913 27081 20947 27115
rect 21189 27081 21223 27115
rect 21557 27081 21591 27115
rect 25237 27081 25271 27115
rect 13369 27013 13403 27047
rect 13461 27013 13495 27047
rect 15853 27013 15887 27047
rect 24317 27013 24351 27047
rect 8309 26945 8343 26979
rect 9413 26945 9447 26979
rect 10517 26945 10551 26979
rect 11897 26945 11931 26979
rect 15117 26945 15151 26979
rect 15209 26945 15243 26979
rect 16313 26945 16347 26979
rect 16865 26945 16899 26979
rect 18061 26945 18095 26979
rect 20269 26945 20303 26979
rect 22017 26945 22051 26979
rect 24593 26945 24627 26979
rect 13553 26877 13587 26911
rect 15393 26877 15427 26911
rect 18337 26877 18371 26911
rect 22293 26877 22327 26911
rect 14749 26809 14783 26843
rect 8953 26741 8987 26775
rect 10057 26741 10091 26775
rect 14381 26741 14415 26775
rect 16129 26741 16163 26775
rect 17509 26741 17543 26775
rect 19809 26741 19843 26775
rect 23765 26741 23799 26775
rect 8585 26537 8619 26571
rect 10517 26537 10551 26571
rect 16313 26537 16347 26571
rect 19704 26537 19738 26571
rect 9137 26469 9171 26503
rect 12081 26469 12115 26503
rect 13553 26469 13587 26503
rect 14105 26469 14139 26503
rect 21189 26469 21223 26503
rect 24593 26469 24627 26503
rect 12633 26401 12667 26435
rect 15025 26401 15059 26435
rect 19441 26401 19475 26435
rect 22293 26401 22327 26435
rect 24041 26401 24075 26435
rect 25237 26401 25271 26435
rect 6837 26333 6871 26367
rect 7941 26333 7975 26367
rect 9229 26333 9263 26367
rect 9873 26333 9907 26367
rect 10977 26333 11011 26367
rect 12449 26333 12483 26367
rect 12541 26333 12575 26367
rect 13737 26333 13771 26367
rect 15669 26333 15703 26367
rect 16773 26333 16807 26367
rect 17969 26333 18003 26367
rect 18981 26333 19015 26367
rect 24961 26333 24995 26367
rect 25053 26333 25087 26367
rect 7481 26265 7515 26299
rect 11621 26265 11655 26299
rect 14841 26265 14875 26299
rect 17417 26265 17451 26299
rect 21649 26265 21683 26299
rect 22569 26265 22603 26299
rect 14473 26197 14507 26231
rect 14933 26197 14967 26231
rect 18613 26197 18647 26231
rect 15393 25993 15427 26027
rect 15485 25993 15519 26027
rect 17233 25993 17267 26027
rect 18429 25993 18463 26027
rect 18521 25993 18555 26027
rect 21281 25993 21315 26027
rect 21557 25993 21591 26027
rect 9689 25925 9723 25959
rect 19073 25925 19107 25959
rect 23397 25925 23431 25959
rect 7205 25857 7239 25891
rect 8309 25857 8343 25891
rect 9413 25857 9447 25891
rect 11713 25857 11747 25891
rect 12817 25857 12851 25891
rect 16129 25857 16163 25891
rect 19533 25857 19567 25891
rect 20177 25857 20211 25891
rect 20637 25857 20671 25891
rect 22017 25857 22051 25891
rect 23121 25857 23155 25891
rect 12357 25789 12391 25823
rect 13093 25789 13127 25823
rect 15577 25789 15611 25823
rect 16313 25789 16347 25823
rect 17325 25789 17359 25823
rect 17417 25789 17451 25823
rect 18705 25789 18739 25823
rect 24869 25789 24903 25823
rect 16405 25721 16439 25755
rect 18061 25721 18095 25755
rect 7849 25653 7883 25687
rect 8953 25653 8987 25687
rect 11161 25653 11195 25687
rect 14565 25653 14599 25687
rect 15025 25653 15059 25687
rect 16865 25653 16899 25687
rect 22661 25653 22695 25687
rect 25237 25653 25271 25687
rect 25421 25653 25455 25687
rect 9394 25449 9428 25483
rect 10885 25449 10919 25483
rect 13553 25449 13587 25483
rect 14473 25449 14507 25483
rect 18705 25449 18739 25483
rect 19073 25449 19107 25483
rect 20177 25449 20211 25483
rect 25237 25449 25271 25483
rect 17601 25381 17635 25415
rect 9137 25313 9171 25347
rect 11345 25313 11379 25347
rect 11621 25313 11655 25347
rect 14933 25313 14967 25347
rect 15025 25313 15059 25347
rect 16221 25313 16255 25347
rect 22017 25313 22051 25347
rect 7941 25245 7975 25279
rect 13737 25245 13771 25279
rect 16129 25245 16163 25279
rect 16957 25245 16991 25279
rect 18061 25245 18095 25279
rect 19533 25245 19567 25279
rect 20729 25245 20763 25279
rect 21925 25245 21959 25279
rect 22661 25245 22695 25279
rect 24593 25245 24627 25279
rect 14841 25177 14875 25211
rect 23857 25177 23891 25211
rect 8585 25109 8619 25143
rect 13093 25109 13127 25143
rect 15669 25109 15703 25143
rect 16037 25109 16071 25143
rect 20821 25109 20855 25143
rect 21465 25109 21499 25143
rect 21833 25109 21867 25143
rect 14473 24905 14507 24939
rect 16405 24905 16439 24939
rect 17233 24905 17267 24939
rect 17325 24905 17359 24939
rect 17877 24905 17911 24939
rect 21833 24905 21867 24939
rect 22753 24905 22787 24939
rect 14381 24837 14415 24871
rect 18889 24837 18923 24871
rect 7481 24769 7515 24803
rect 8585 24769 8619 24803
rect 11713 24769 11747 24803
rect 13185 24769 13219 24803
rect 13277 24769 13311 24803
rect 15209 24769 15243 24803
rect 15853 24769 15887 24803
rect 19717 24769 19751 24803
rect 8125 24701 8159 24735
rect 8861 24701 8895 24735
rect 10977 24701 11011 24735
rect 13369 24701 13403 24735
rect 14657 24701 14691 24735
rect 17417 24701 17451 24735
rect 18153 24701 18187 24735
rect 18981 24701 19015 24735
rect 19073 24701 19107 24735
rect 19993 24701 20027 24735
rect 22845 24701 22879 24735
rect 22937 24701 22971 24735
rect 23581 24701 23615 24735
rect 23857 24701 23891 24735
rect 18521 24633 18555 24667
rect 10333 24565 10367 24599
rect 12357 24565 12391 24599
rect 12817 24565 12851 24599
rect 14013 24565 14047 24599
rect 16221 24565 16255 24599
rect 16865 24565 16899 24599
rect 21465 24565 21499 24599
rect 22109 24565 22143 24599
rect 22385 24565 22419 24599
rect 25329 24565 25363 24599
rect 10057 24361 10091 24395
rect 15301 24361 15335 24395
rect 21557 24361 21591 24395
rect 25237 24361 25271 24395
rect 14933 24293 14967 24327
rect 10701 24225 10735 24259
rect 11529 24225 11563 24259
rect 18705 24225 18739 24259
rect 20085 24225 20119 24259
rect 5733 24157 5767 24191
rect 6837 24157 6871 24191
rect 7941 24157 7975 24191
rect 10425 24157 10459 24191
rect 11253 24157 11287 24191
rect 14289 24157 14323 24191
rect 15485 24157 15519 24191
rect 19809 24157 19843 24191
rect 20913 24157 20947 24191
rect 22017 24157 22051 24191
rect 24593 24157 24627 24191
rect 8585 24089 8619 24123
rect 9413 24089 9447 24123
rect 15945 24089 15979 24123
rect 20453 24089 20487 24123
rect 22293 24089 22327 24123
rect 6377 24021 6411 24055
rect 7481 24021 7515 24055
rect 10517 24021 10551 24055
rect 13001 24021 13035 24055
rect 13553 24021 13587 24055
rect 15669 24021 15703 24055
rect 17233 24021 17267 24055
rect 18153 24021 18187 24055
rect 18521 24021 18555 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 19901 24021 19935 24055
rect 23765 24021 23799 24055
rect 24041 24021 24075 24055
rect 6469 23817 6503 23851
rect 9137 23817 9171 23851
rect 9597 23817 9631 23851
rect 11161 23817 11195 23851
rect 11805 23817 11839 23851
rect 13093 23817 13127 23851
rect 13921 23817 13955 23851
rect 15853 23817 15887 23851
rect 21833 23817 21867 23851
rect 22385 23817 22419 23851
rect 22477 23817 22511 23851
rect 24961 23817 24995 23851
rect 14013 23749 14047 23783
rect 19349 23749 19383 23783
rect 25329 23749 25363 23783
rect 25513 23749 25547 23783
rect 6929 23681 6963 23715
rect 9505 23681 9539 23715
rect 10517 23681 10551 23715
rect 11989 23681 12023 23715
rect 12449 23681 12483 23715
rect 14749 23681 14783 23715
rect 16865 23681 16899 23715
rect 17969 23681 18003 23715
rect 19073 23681 19107 23715
rect 21465 23681 21499 23715
rect 7205 23613 7239 23647
rect 9689 23613 9723 23647
rect 14197 23613 14231 23647
rect 20821 23613 20855 23647
rect 22661 23613 22695 23647
rect 23213 23613 23247 23647
rect 23489 23613 23523 23647
rect 8309 23477 8343 23511
rect 13553 23477 13587 23511
rect 15393 23477 15427 23511
rect 17509 23477 17543 23511
rect 18613 23477 18647 23511
rect 21281 23477 21315 23511
rect 22017 23477 22051 23511
rect 8585 23273 8619 23307
rect 13001 23273 13035 23307
rect 22293 23273 22327 23307
rect 7205 23205 7239 23239
rect 18889 23205 18923 23239
rect 6009 23137 6043 23171
rect 9137 23137 9171 23171
rect 12265 23137 12299 23171
rect 13553 23137 13587 23171
rect 14565 23137 14599 23171
rect 17049 23137 17083 23171
rect 17785 23137 17819 23171
rect 19349 23137 19383 23171
rect 20545 23137 20579 23171
rect 22109 23137 22143 23171
rect 23857 23137 23891 23171
rect 25145 23137 25179 23171
rect 6285 23069 6319 23103
rect 7297 23069 7331 23103
rect 7941 23069 7975 23103
rect 12081 23069 12115 23103
rect 12173 23069 12207 23103
rect 14289 23069 14323 23103
rect 16957 23069 16991 23103
rect 18245 23069 18279 23103
rect 20269 23069 20303 23103
rect 21097 23069 21131 23103
rect 22661 23069 22695 23103
rect 25053 23069 25087 23103
rect 9413 23001 9447 23035
rect 13369 23001 13403 23035
rect 20361 23001 20395 23035
rect 24961 23001 24995 23035
rect 10885 22933 10919 22967
rect 11713 22933 11747 22967
rect 13461 22933 13495 22967
rect 16037 22933 16071 22967
rect 16497 22933 16531 22967
rect 16865 22933 16899 22967
rect 17601 22933 17635 22967
rect 17969 22933 18003 22967
rect 19533 22933 19567 22967
rect 19901 22933 19935 22967
rect 21741 22933 21775 22967
rect 24593 22933 24627 22967
rect 12081 22729 12115 22763
rect 15761 22729 15795 22763
rect 17509 22729 17543 22763
rect 18429 22729 18463 22763
rect 19165 22729 19199 22763
rect 19901 22729 19935 22763
rect 19993 22729 20027 22763
rect 21373 22729 21407 22763
rect 6653 22661 6687 22695
rect 12173 22661 12207 22695
rect 18337 22661 18371 22695
rect 18981 22661 19015 22695
rect 8585 22593 8619 22627
rect 12909 22593 12943 22627
rect 16865 22593 16899 22627
rect 20729 22593 20763 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 7297 22525 7331 22559
rect 7573 22525 7607 22559
rect 8861 22525 8895 22559
rect 10977 22525 11011 22559
rect 12265 22525 12299 22559
rect 14013 22525 14047 22559
rect 14289 22525 14323 22559
rect 16405 22525 16439 22559
rect 18521 22525 18555 22559
rect 20085 22525 20119 22559
rect 23305 22525 23339 22559
rect 24777 22525 24811 22559
rect 7205 22457 7239 22491
rect 10333 22389 10367 22423
rect 10701 22389 10735 22423
rect 11713 22389 11747 22423
rect 13553 22389 13587 22423
rect 17969 22389 18003 22423
rect 19533 22389 19567 22423
rect 19257 22185 19291 22219
rect 21005 22185 21039 22219
rect 21728 22185 21762 22219
rect 6837 22049 6871 22083
rect 8585 22049 8619 22083
rect 10793 22049 10827 22083
rect 15301 22049 15335 22083
rect 16497 22049 16531 22083
rect 19441 22049 19475 22083
rect 20453 22049 20487 22083
rect 21465 22049 21499 22083
rect 25053 22049 25087 22083
rect 25237 22049 25271 22083
rect 6377 21981 6411 22015
rect 9137 21981 9171 22015
rect 10701 21981 10735 22015
rect 11989 21981 12023 22015
rect 13093 21981 13127 22015
rect 15117 21981 15151 22015
rect 16313 21981 16347 22015
rect 16405 21981 16439 22015
rect 17141 21981 17175 22015
rect 18245 21981 18279 22015
rect 20177 21981 20211 22015
rect 20269 21981 20303 22015
rect 23949 21981 23983 22015
rect 7113 21913 7147 21947
rect 6193 21845 6227 21879
rect 9781 21845 9815 21879
rect 10241 21845 10275 21879
rect 10609 21845 10643 21879
rect 11529 21845 11563 21879
rect 12633 21845 12667 21879
rect 13737 21845 13771 21879
rect 14749 21845 14783 21879
rect 15209 21845 15243 21879
rect 15945 21845 15979 21879
rect 17785 21845 17819 21879
rect 18889 21845 18923 21879
rect 19809 21845 19843 21879
rect 21097 21845 21131 21879
rect 23213 21845 23247 21879
rect 23765 21845 23799 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 8585 21641 8619 21675
rect 9965 21641 9999 21675
rect 10425 21641 10459 21675
rect 10885 21641 10919 21675
rect 15761 21641 15795 21675
rect 19809 21641 19843 21675
rect 25421 21641 25455 21675
rect 13185 21573 13219 21607
rect 16037 21573 16071 21607
rect 19165 21573 19199 21607
rect 22385 21573 22419 21607
rect 22477 21573 22511 21607
rect 25329 21573 25363 21607
rect 5457 21505 5491 21539
rect 6837 21505 6871 21539
rect 7941 21505 7975 21539
rect 9321 21505 9355 21539
rect 10793 21505 10827 21539
rect 12081 21505 12115 21539
rect 15117 21505 15151 21539
rect 16865 21505 16899 21539
rect 20269 21505 20303 21539
rect 5181 21437 5215 21471
rect 10977 21437 11011 21471
rect 12173 21437 12207 21471
rect 12265 21437 12299 21471
rect 12909 21437 12943 21471
rect 17141 21437 17175 21471
rect 21281 21437 21315 21471
rect 22569 21437 22603 21471
rect 23213 21437 23247 21471
rect 23489 21437 23523 21471
rect 6469 21369 6503 21403
rect 7481 21301 7515 21335
rect 11713 21301 11747 21335
rect 14657 21301 14691 21335
rect 16313 21301 16347 21335
rect 16497 21301 16531 21335
rect 18613 21301 18647 21335
rect 19257 21301 19291 21335
rect 22017 21301 22051 21335
rect 24961 21301 24995 21335
rect 10425 21097 10459 21131
rect 13921 21029 13955 21063
rect 15301 21029 15335 21063
rect 16405 21029 16439 21063
rect 18613 21029 18647 21063
rect 18981 21029 19015 21063
rect 19441 21029 19475 21063
rect 21833 21029 21867 21063
rect 22293 21029 22327 21063
rect 24593 21029 24627 21063
rect 8585 20961 8619 20995
rect 10977 20961 11011 20995
rect 11621 20961 11655 20995
rect 20085 20961 20119 20995
rect 21281 20961 21315 20995
rect 23857 20961 23891 20995
rect 25145 20961 25179 20995
rect 5733 20893 5767 20927
rect 6837 20893 6871 20927
rect 7941 20893 7975 20927
rect 9321 20893 9355 20927
rect 9965 20893 9999 20927
rect 14657 20893 14691 20927
rect 15761 20893 15795 20927
rect 16865 20893 16899 20927
rect 17509 20893 17543 20927
rect 17969 20893 18003 20927
rect 19901 20893 19935 20927
rect 22017 20893 22051 20927
rect 22845 20893 22879 20927
rect 10793 20825 10827 20859
rect 11897 20825 11931 20859
rect 21097 20825 21131 20859
rect 25053 20825 25087 20859
rect 5089 20757 5123 20791
rect 6377 20757 6411 20791
rect 7481 20757 7515 20791
rect 10885 20757 10919 20791
rect 13369 20757 13403 20791
rect 13645 20757 13679 20791
rect 14197 20757 14231 20791
rect 14381 20757 14415 20791
rect 19809 20757 19843 20791
rect 20637 20757 20671 20791
rect 21005 20757 21039 20791
rect 24961 20757 24995 20791
rect 6009 20553 6043 20587
rect 10793 20553 10827 20587
rect 12357 20553 12391 20587
rect 19165 20553 19199 20587
rect 19349 20553 19383 20587
rect 21465 20553 21499 20587
rect 21833 20553 21867 20587
rect 22477 20553 22511 20587
rect 23213 20553 23247 20587
rect 25329 20553 25363 20587
rect 4905 20485 4939 20519
rect 5365 20417 5399 20451
rect 6837 20417 6871 20451
rect 8217 20417 8251 20451
rect 11713 20417 11747 20451
rect 12817 20417 12851 20451
rect 14105 20417 14139 20451
rect 16957 20417 16991 20451
rect 19993 20417 20027 20451
rect 20821 20417 20855 20451
rect 22385 20417 22419 20451
rect 23581 20417 23615 20451
rect 4353 20349 4387 20383
rect 7481 20349 7515 20383
rect 8493 20349 8527 20383
rect 10241 20349 10275 20383
rect 14565 20349 14599 20383
rect 14841 20349 14875 20383
rect 17233 20349 17267 20383
rect 20085 20349 20119 20383
rect 20269 20349 20303 20383
rect 22661 20349 22695 20383
rect 23857 20349 23891 20383
rect 22017 20281 22051 20315
rect 13461 20213 13495 20247
rect 13921 20213 13955 20247
rect 16313 20213 16347 20247
rect 18705 20213 18739 20247
rect 19625 20213 19659 20247
rect 23121 20213 23155 20247
rect 7849 20009 7883 20043
rect 9946 20009 9980 20043
rect 13645 20009 13679 20043
rect 17049 20009 17083 20043
rect 18797 20009 18831 20043
rect 19073 20009 19107 20043
rect 25237 20009 25271 20043
rect 6285 19941 6319 19975
rect 4353 19873 4387 19907
rect 7389 19873 7423 19907
rect 8401 19873 8435 19907
rect 14473 19873 14507 19907
rect 15761 19873 15795 19907
rect 18245 19873 18279 19907
rect 23857 19873 23891 19907
rect 4629 19805 4663 19839
rect 5641 19805 5675 19839
rect 6745 19805 6779 19839
rect 9689 19805 9723 19839
rect 12173 19805 12207 19839
rect 12633 19805 12667 19839
rect 13921 19805 13955 19839
rect 14289 19805 14323 19839
rect 16405 19805 16439 19839
rect 18061 19805 18095 19839
rect 19441 19805 19475 19839
rect 20821 19805 20855 19839
rect 22661 19805 22695 19839
rect 24593 19805 24627 19839
rect 8217 19737 8251 19771
rect 15669 19737 15703 19771
rect 18705 19737 18739 19771
rect 22017 19737 22051 19771
rect 8309 19669 8343 19703
rect 11437 19669 11471 19703
rect 11989 19669 12023 19703
rect 13277 19669 13311 19703
rect 15209 19669 15243 19703
rect 15577 19669 15611 19703
rect 17601 19669 17635 19703
rect 17969 19669 18003 19703
rect 20085 19669 20119 19703
rect 20361 19669 20395 19703
rect 4997 19465 5031 19499
rect 6009 19465 6043 19499
rect 6653 19465 6687 19499
rect 9045 19465 9079 19499
rect 9597 19465 9631 19499
rect 10977 19465 11011 19499
rect 12265 19465 12299 19499
rect 15853 19465 15887 19499
rect 17509 19465 17543 19499
rect 17969 19465 18003 19499
rect 24225 19465 24259 19499
rect 24685 19465 24719 19499
rect 25513 19465 25547 19499
rect 10057 19397 10091 19431
rect 3985 19329 4019 19363
rect 5365 19329 5399 19363
rect 7297 19329 7331 19363
rect 9965 19329 9999 19363
rect 11161 19329 11195 19363
rect 12633 19329 12667 19363
rect 12725 19329 12759 19363
rect 14105 19329 14139 19363
rect 16865 19329 16899 19363
rect 18153 19329 18187 19363
rect 18613 19329 18647 19363
rect 19717 19329 19751 19363
rect 22017 19329 22051 19363
rect 24593 19329 24627 19363
rect 3709 19261 3743 19295
rect 4813 19261 4847 19295
rect 7573 19261 7607 19295
rect 10241 19261 10275 19295
rect 12817 19261 12851 19295
rect 13461 19261 13495 19295
rect 14381 19261 14415 19295
rect 19993 19261 20027 19295
rect 22293 19261 22327 19295
rect 23765 19261 23799 19295
rect 24777 19261 24811 19295
rect 25237 19261 25271 19295
rect 24041 19193 24075 19227
rect 10609 19125 10643 19159
rect 11529 19125 11563 19159
rect 11805 19125 11839 19159
rect 11989 19125 12023 19159
rect 16221 19125 16255 19159
rect 16405 19125 16439 19159
rect 19257 19125 19291 19159
rect 21465 19125 21499 19159
rect 21465 18921 21499 18955
rect 21925 18921 21959 18955
rect 25237 18921 25271 18955
rect 6009 18853 6043 18887
rect 9597 18853 9631 18887
rect 10793 18853 10827 18887
rect 18153 18853 18187 18887
rect 18889 18853 18923 18887
rect 6653 18785 6687 18819
rect 8401 18785 8435 18819
rect 10149 18785 10183 18819
rect 11253 18785 11287 18819
rect 11437 18785 11471 18819
rect 11989 18785 12023 18819
rect 16497 18785 16531 18819
rect 16589 18785 16623 18819
rect 20821 18785 20855 18819
rect 22293 18785 22327 18819
rect 4261 18717 4295 18751
rect 4905 18717 4939 18751
rect 5365 18717 5399 18751
rect 9965 18717 9999 18751
rect 10057 18717 10091 18751
rect 14289 18717 14323 18751
rect 15577 18717 15611 18751
rect 16405 18717 16439 18751
rect 17233 18717 17267 18751
rect 19533 18717 19567 18751
rect 20545 18717 20579 18751
rect 21649 18717 21683 18751
rect 24593 18717 24627 18751
rect 3157 18649 3191 18683
rect 3249 18649 3283 18683
rect 6929 18649 6963 18683
rect 12265 18649 12299 18683
rect 18705 18649 18739 18683
rect 19717 18649 19751 18683
rect 22569 18649 22603 18683
rect 4077 18581 4111 18615
rect 4721 18581 4755 18615
rect 9045 18581 9079 18615
rect 9229 18581 9263 18615
rect 11161 18581 11195 18615
rect 13737 18581 13771 18615
rect 14933 18581 14967 18615
rect 15393 18581 15427 18615
rect 16037 18581 16071 18615
rect 17877 18581 17911 18615
rect 20177 18581 20211 18615
rect 20637 18581 20671 18615
rect 24041 18581 24075 18615
rect 6009 18377 6043 18411
rect 9781 18377 9815 18411
rect 10425 18377 10459 18411
rect 12357 18377 12391 18411
rect 12909 18377 12943 18411
rect 13277 18377 13311 18411
rect 15209 18377 15243 18411
rect 19717 18377 19751 18411
rect 20177 18377 20211 18411
rect 21465 18377 21499 18411
rect 4537 18309 4571 18343
rect 10057 18309 10091 18343
rect 10793 18309 10827 18343
rect 10885 18309 10919 18343
rect 16313 18309 16347 18343
rect 17141 18309 17175 18343
rect 3985 18241 4019 18275
rect 5365 18241 5399 18275
rect 6929 18241 6963 18275
rect 8033 18241 8067 18275
rect 11713 18241 11747 18275
rect 14565 18241 14599 18275
rect 15669 18241 15703 18275
rect 16865 18241 16899 18275
rect 19073 18241 19107 18275
rect 20821 18241 20855 18275
rect 22017 18241 22051 18275
rect 23489 18241 23523 18275
rect 4721 18173 4755 18207
rect 7573 18173 7607 18207
rect 8309 18173 8343 18207
rect 11069 18173 11103 18207
rect 13369 18173 13403 18207
rect 13461 18173 13495 18207
rect 22661 18173 22695 18207
rect 23765 18173 23799 18207
rect 3801 18037 3835 18071
rect 13921 18037 13955 18071
rect 14197 18037 14231 18071
rect 18613 18037 18647 18071
rect 23029 18037 23063 18071
rect 25237 18037 25271 18071
rect 9137 17833 9171 17867
rect 13001 17833 13035 17867
rect 15301 17833 15335 17867
rect 15761 17833 15795 17867
rect 21097 17833 21131 17867
rect 22201 17833 22235 17867
rect 5181 17765 5215 17799
rect 3249 17697 3283 17731
rect 4261 17697 4295 17731
rect 5825 17697 5859 17731
rect 6469 17697 6503 17731
rect 9689 17697 9723 17731
rect 10793 17697 10827 17731
rect 13553 17697 13587 17731
rect 17417 17697 17451 17731
rect 18613 17697 18647 17731
rect 20085 17697 20119 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 4721 17629 4755 17663
rect 5365 17629 5399 17663
rect 6837 17629 6871 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 10517 17629 10551 17663
rect 13369 17629 13403 17663
rect 14105 17629 14139 17663
rect 14657 17629 14691 17663
rect 16129 17629 16163 17663
rect 17141 17629 17175 17663
rect 18521 17629 18555 17663
rect 19533 17629 19567 17663
rect 20453 17629 20487 17663
rect 21557 17629 21591 17663
rect 22661 17629 22695 17663
rect 6377 17561 6411 17595
rect 9505 17561 9539 17595
rect 9597 17561 9631 17595
rect 10149 17561 10183 17595
rect 12541 17561 12575 17595
rect 13461 17561 13495 17595
rect 14289 17561 14323 17595
rect 16313 17561 16347 17595
rect 4537 17493 4571 17527
rect 7481 17493 7515 17527
rect 16773 17493 16807 17527
rect 17233 17493 17267 17527
rect 18061 17493 18095 17527
rect 18429 17493 18463 17527
rect 19625 17493 19659 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 6009 17289 6043 17323
rect 6377 17289 6411 17323
rect 8677 17289 8711 17323
rect 9965 17289 9999 17323
rect 10425 17289 10459 17323
rect 10885 17289 10919 17323
rect 13829 17289 13863 17323
rect 18889 17289 18923 17323
rect 20361 17289 20395 17323
rect 22937 17289 22971 17323
rect 23581 17289 23615 17323
rect 9045 17221 9079 17255
rect 10149 17221 10183 17255
rect 13185 17221 13219 17255
rect 14197 17221 14231 17255
rect 16129 17221 16163 17255
rect 3617 17153 3651 17187
rect 4077 17153 4111 17187
rect 5365 17153 5399 17187
rect 7573 17153 7607 17187
rect 10793 17153 10827 17187
rect 12449 17153 12483 17187
rect 15025 17153 15059 17187
rect 17417 17153 17451 17187
rect 18245 17153 18279 17187
rect 19717 17153 19751 17187
rect 20821 17153 20855 17187
rect 21465 17153 21499 17187
rect 22109 17153 22143 17187
rect 22845 17153 22879 17187
rect 23949 17153 23983 17187
rect 2789 17085 2823 17119
rect 4353 17085 4387 17119
rect 6561 17085 6595 17119
rect 6929 17085 6963 17119
rect 9137 17085 9171 17119
rect 9321 17085 9355 17119
rect 10977 17085 11011 17119
rect 11805 17085 11839 17119
rect 14289 17085 14323 17119
rect 14473 17085 14507 17119
rect 17509 17085 17543 17119
rect 17693 17085 17727 17119
rect 21925 17085 21959 17119
rect 23121 17085 23155 17119
rect 24777 17085 24811 17119
rect 15669 17017 15703 17051
rect 19349 17017 19383 17051
rect 22477 17017 22511 17051
rect 3433 16949 3467 16983
rect 8217 16949 8251 16983
rect 9781 16949 9815 16983
rect 16681 16949 16715 16983
rect 17049 16949 17083 16983
rect 19165 16949 19199 16983
rect 8125 16745 8159 16779
rect 14197 16745 14231 16779
rect 17417 16745 17451 16779
rect 19349 16745 19383 16779
rect 21005 16745 21039 16779
rect 22201 16745 22235 16779
rect 8677 16677 8711 16711
rect 16405 16677 16439 16711
rect 17141 16677 17175 16711
rect 3985 16609 4019 16643
rect 4261 16609 4295 16643
rect 6653 16609 6687 16643
rect 9597 16609 9631 16643
rect 9689 16609 9723 16643
rect 11253 16609 11287 16643
rect 13277 16609 13311 16643
rect 14657 16609 14691 16643
rect 18521 16609 18555 16643
rect 18981 16609 19015 16643
rect 20545 16609 20579 16643
rect 5273 16541 5307 16575
rect 5917 16541 5951 16575
rect 6377 16541 6411 16575
rect 10517 16541 10551 16575
rect 11805 16541 11839 16575
rect 12265 16541 12299 16575
rect 17785 16541 17819 16575
rect 19717 16541 19751 16575
rect 21557 16541 21591 16575
rect 22661 16541 22695 16575
rect 24593 16541 24627 16575
rect 25237 16541 25271 16575
rect 14933 16473 14967 16507
rect 16957 16473 16991 16507
rect 23857 16473 23891 16507
rect 3249 16405 3283 16439
rect 8493 16405 8527 16439
rect 9137 16405 9171 16439
rect 9505 16405 9539 16439
rect 10149 16405 10183 16439
rect 12081 16405 12115 16439
rect 12725 16405 12759 16439
rect 13093 16405 13127 16439
rect 13185 16405 13219 16439
rect 13829 16405 13863 16439
rect 14381 16405 14415 16439
rect 16681 16405 16715 16439
rect 21281 16405 21315 16439
rect 6469 16201 6503 16235
rect 10425 16201 10459 16235
rect 10885 16201 10919 16235
rect 13921 16201 13955 16235
rect 14289 16201 14323 16235
rect 15669 16201 15703 16235
rect 18061 16201 18095 16235
rect 21189 16201 21223 16235
rect 4077 16133 4111 16167
rect 4261 16133 4295 16167
rect 8217 16133 8251 16167
rect 10793 16133 10827 16167
rect 17509 16133 17543 16167
rect 25145 16133 25179 16167
rect 3617 16065 3651 16099
rect 4905 16065 4939 16099
rect 5365 16065 5399 16099
rect 6848 16065 6882 16099
rect 7941 16065 7975 16099
rect 16313 16065 16347 16099
rect 16865 16065 16899 16099
rect 18429 16065 18463 16099
rect 21097 16065 21131 16099
rect 22109 16065 22143 16099
rect 23949 16065 23983 16099
rect 3433 15997 3467 16031
rect 9965 15997 9999 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 14381 15997 14415 16031
rect 14473 15997 14507 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 17969 15997 18003 16031
rect 18705 15997 18739 16031
rect 21373 15997 21407 16031
rect 23305 15997 23339 16031
rect 1593 15929 1627 15963
rect 15301 15929 15335 15963
rect 20729 15929 20763 15963
rect 2237 15861 2271 15895
rect 4721 15861 4755 15895
rect 6009 15861 6043 15895
rect 7481 15861 7515 15895
rect 13461 15861 13495 15895
rect 15025 15861 15059 15895
rect 20177 15861 20211 15895
rect 3341 15657 3375 15691
rect 5089 15657 5123 15691
rect 6193 15657 6227 15691
rect 8769 15657 8803 15691
rect 9137 15657 9171 15691
rect 11805 15657 11839 15691
rect 2881 15589 2915 15623
rect 8401 15589 8435 15623
rect 9781 15589 9815 15623
rect 11345 15589 11379 15623
rect 1961 15521 1995 15555
rect 6653 15521 6687 15555
rect 10333 15521 10367 15555
rect 12357 15521 12391 15555
rect 13645 15521 13679 15555
rect 14841 15521 14875 15555
rect 16313 15521 16347 15555
rect 16589 15521 16623 15555
rect 20361 15521 20395 15555
rect 22109 15521 22143 15555
rect 2605 15453 2639 15487
rect 4445 15453 4479 15487
rect 5549 15453 5583 15487
rect 9321 15453 9355 15487
rect 10149 15453 10183 15487
rect 13369 15453 13403 15487
rect 14657 15453 14691 15487
rect 15577 15453 15611 15487
rect 18613 15453 18647 15487
rect 19993 15453 20027 15487
rect 22661 15453 22695 15487
rect 24685 15453 24719 15487
rect 1685 15385 1719 15419
rect 3249 15385 3283 15419
rect 4169 15385 4203 15419
rect 6929 15385 6963 15419
rect 11161 15385 11195 15419
rect 14749 15385 14783 15419
rect 15761 15385 15795 15419
rect 18797 15385 18831 15419
rect 19533 15385 19567 15419
rect 19717 15385 19751 15419
rect 20637 15385 20671 15419
rect 23857 15385 23891 15419
rect 1501 15317 1535 15351
rect 2053 15317 2087 15351
rect 2237 15317 2271 15351
rect 2421 15317 2455 15351
rect 2973 15317 3007 15351
rect 3617 15317 3651 15351
rect 3893 15317 3927 15351
rect 10241 15317 10275 15351
rect 12173 15317 12207 15351
rect 12265 15317 12299 15351
rect 13001 15317 13035 15351
rect 13461 15317 13495 15351
rect 14289 15317 14323 15351
rect 18061 15317 18095 15351
rect 25329 15317 25363 15351
rect 4905 15113 4939 15147
rect 14197 15113 14231 15147
rect 15393 15113 15427 15147
rect 16313 15113 16347 15147
rect 16865 15113 16899 15147
rect 24041 15113 24075 15147
rect 10057 15045 10091 15079
rect 17233 15045 17267 15079
rect 21373 15045 21407 15079
rect 3249 14977 3283 15011
rect 4261 14977 4295 15011
rect 5365 14977 5399 15011
rect 6929 14977 6963 15011
rect 8033 14977 8067 15011
rect 10517 14977 10551 15011
rect 11161 14977 11195 15011
rect 11713 14977 11747 15011
rect 12817 14977 12851 15011
rect 13553 14977 13587 15011
rect 14565 14977 14599 15011
rect 15669 14977 15703 15011
rect 17877 14977 17911 15011
rect 18245 14977 18279 15011
rect 19349 14977 19383 15011
rect 24409 14977 24443 15011
rect 24685 14977 24719 15011
rect 1961 14909 1995 14943
rect 8309 14909 8343 14943
rect 14657 14909 14691 14943
rect 14841 14909 14875 14943
rect 17325 14909 17359 14943
rect 17509 14909 17543 14943
rect 19625 14909 19659 14943
rect 22017 14909 22051 14943
rect 22293 14909 22327 14943
rect 2421 14841 2455 14875
rect 6009 14841 6043 14875
rect 6469 14841 6503 14875
rect 6653 14841 6687 14875
rect 1501 14773 1535 14807
rect 1685 14773 1719 14807
rect 1869 14773 1903 14807
rect 2145 14773 2179 14807
rect 2605 14773 2639 14807
rect 2881 14773 2915 14807
rect 3801 14773 3835 14807
rect 7573 14773 7607 14807
rect 12357 14773 12391 14807
rect 18889 14773 18923 14807
rect 21097 14773 21131 14807
rect 21557 14773 21591 14807
rect 23765 14773 23799 14807
rect 3893 14569 3927 14603
rect 6377 14569 6411 14603
rect 10406 14569 10440 14603
rect 12633 14569 12667 14603
rect 15485 14569 15519 14603
rect 16589 14569 16623 14603
rect 20637 14569 20671 14603
rect 23949 14569 23983 14603
rect 3249 14501 3283 14535
rect 8585 14501 8619 14535
rect 14197 14501 14231 14535
rect 9229 14433 9263 14467
rect 9505 14433 9539 14467
rect 10149 14433 10183 14467
rect 12173 14433 12207 14467
rect 13277 14433 13311 14467
rect 13921 14433 13955 14467
rect 20085 14433 20119 14467
rect 21281 14433 21315 14467
rect 21649 14433 21683 14467
rect 22201 14433 22235 14467
rect 2053 14365 2087 14399
rect 2605 14365 2639 14399
rect 3433 14365 3467 14399
rect 3985 14365 4019 14399
rect 4721 14365 4755 14399
rect 5733 14365 5767 14399
rect 6837 14365 6871 14399
rect 7975 14365 8009 14399
rect 14473 14365 14507 14399
rect 15945 14365 15979 14399
rect 17049 14365 17083 14399
rect 18245 14365 18279 14399
rect 19533 14365 19567 14399
rect 21097 14365 21131 14399
rect 21833 14365 21867 14399
rect 24593 14365 24627 14399
rect 2789 14297 2823 14331
rect 5273 14297 5307 14331
rect 13001 14297 13035 14331
rect 13093 14297 13127 14331
rect 15577 14297 15611 14331
rect 22477 14297 22511 14331
rect 1501 14229 1535 14263
rect 1869 14229 1903 14263
rect 7481 14229 7515 14263
rect 8953 14229 8987 14263
rect 13645 14229 13679 14263
rect 15117 14229 15151 14263
rect 17693 14229 17727 14263
rect 18889 14229 18923 14263
rect 21005 14229 21039 14263
rect 25237 14229 25271 14263
rect 1685 14025 1719 14059
rect 6009 14025 6043 14059
rect 6469 14025 6503 14059
rect 9597 14025 9631 14059
rect 10425 14025 10459 14059
rect 10885 14025 10919 14059
rect 12357 14025 12391 14059
rect 12817 14025 12851 14059
rect 13185 14025 13219 14059
rect 13277 14025 13311 14059
rect 16865 14025 16899 14059
rect 17233 14025 17267 14059
rect 17969 14025 18003 14059
rect 19073 14025 19107 14059
rect 19349 14025 19383 14059
rect 20177 14025 20211 14059
rect 21281 14025 21315 14059
rect 25053 14025 25087 14059
rect 4905 13957 4939 13991
rect 14289 13957 14323 13991
rect 17325 13957 17359 13991
rect 20821 13957 20855 13991
rect 22109 13957 22143 13991
rect 2329 13889 2363 13923
rect 4261 13889 4295 13923
rect 5365 13889 5399 13923
rect 6745 13889 6779 13923
rect 8953 13889 8987 13923
rect 10793 13889 10827 13923
rect 11713 13889 11747 13923
rect 16405 13889 16439 13923
rect 18061 13889 18095 13923
rect 18429 13889 18463 13923
rect 20085 13889 20119 13923
rect 21097 13889 21131 13923
rect 21465 13889 21499 13923
rect 25237 13889 25271 13923
rect 2605 13821 2639 13855
rect 3617 13821 3651 13855
rect 8493 13821 8527 13855
rect 9689 13821 9723 13855
rect 9781 13821 9815 13855
rect 10977 13821 11011 13855
rect 13369 13821 13403 13855
rect 14013 13821 14047 13855
rect 15761 13821 15795 13855
rect 16037 13821 16071 13855
rect 17417 13821 17451 13855
rect 20269 13821 20303 13855
rect 20913 13821 20947 13855
rect 22845 13821 22879 13855
rect 24593 13821 24627 13855
rect 9229 13753 9263 13787
rect 19717 13753 19751 13787
rect 22293 13753 22327 13787
rect 7008 13685 7042 13719
rect 16221 13685 16255 13719
rect 23108 13685 23142 13719
rect 4077 13481 4111 13515
rect 6285 13481 6319 13515
rect 9137 13481 9171 13515
rect 10425 13481 10459 13515
rect 14197 13481 14231 13515
rect 17601 13481 17635 13515
rect 18889 13481 18923 13515
rect 19349 13481 19383 13515
rect 19441 13481 19475 13515
rect 22109 13481 22143 13515
rect 25237 13481 25271 13515
rect 7389 13413 7423 13447
rect 14841 13413 14875 13447
rect 2513 13345 2547 13379
rect 3249 13345 3283 13379
rect 8309 13345 8343 13379
rect 8401 13345 8435 13379
rect 9689 13345 9723 13379
rect 10977 13345 11011 13379
rect 11529 13345 11563 13379
rect 12265 13345 12299 13379
rect 12357 13345 12391 13379
rect 13645 13345 13679 13379
rect 15853 13345 15887 13379
rect 19993 13345 20027 13379
rect 21281 13345 21315 13379
rect 23857 13345 23891 13379
rect 1777 13277 1811 13311
rect 2329 13277 2363 13311
rect 3065 13277 3099 13311
rect 4261 13277 4295 13311
rect 4537 13277 4571 13311
rect 5641 13277 5675 13311
rect 6745 13277 6779 13311
rect 9505 13277 9539 13311
rect 10793 13277 10827 13311
rect 13461 13277 13495 13311
rect 16497 13277 16531 13311
rect 17785 13277 17819 13311
rect 18245 13277 18279 13311
rect 19901 13277 19935 13311
rect 21189 13277 21223 13311
rect 22017 13277 22051 13311
rect 22661 13277 22695 13311
rect 24593 13277 24627 13311
rect 3801 13209 3835 13243
rect 5181 13209 5215 13243
rect 8217 13209 8251 13243
rect 9597 13209 9631 13243
rect 12173 13209 12207 13243
rect 14657 13209 14691 13243
rect 15669 13209 15703 13243
rect 1593 13141 1627 13175
rect 3617 13141 3651 13175
rect 7849 13141 7883 13175
rect 10885 13141 10919 13175
rect 11805 13141 11839 13175
rect 13001 13141 13035 13175
rect 13369 13141 13403 13175
rect 15301 13141 15335 13175
rect 15761 13141 15795 13175
rect 17141 13141 17175 13175
rect 19809 13141 19843 13175
rect 20729 13141 20763 13175
rect 21097 13141 21131 13175
rect 2605 12937 2639 12971
rect 3893 12937 3927 12971
rect 13093 12937 13127 12971
rect 13461 12937 13495 12971
rect 19257 12937 19291 12971
rect 25237 12937 25271 12971
rect 3249 12869 3283 12903
rect 7481 12869 7515 12903
rect 11713 12869 11747 12903
rect 12449 12869 12483 12903
rect 15945 12869 15979 12903
rect 19073 12869 19107 12903
rect 19625 12869 19659 12903
rect 21097 12869 21131 12903
rect 21649 12869 21683 12903
rect 23305 12869 23339 12903
rect 25053 12869 25087 12903
rect 2145 12801 2179 12835
rect 2789 12801 2823 12835
rect 4261 12801 4295 12835
rect 5365 12801 5399 12835
rect 8309 12801 8343 12835
rect 9413 12801 9447 12835
rect 14749 12801 14783 12835
rect 16037 12801 16071 12835
rect 22109 12801 22143 12835
rect 25421 12801 25455 12835
rect 6837 12733 6871 12767
rect 7573 12733 7607 12767
rect 7665 12733 7699 12767
rect 8953 12733 8987 12767
rect 9689 12733 9723 12767
rect 13553 12733 13587 12767
rect 13737 12733 13771 12767
rect 14841 12733 14875 12767
rect 14933 12733 14967 12767
rect 16129 12733 16163 12767
rect 16865 12733 16899 12767
rect 17141 12733 17175 12767
rect 20453 12733 20487 12767
rect 22293 12733 22327 12767
rect 23029 12733 23063 12767
rect 1685 12665 1719 12699
rect 1961 12665 1995 12699
rect 6469 12665 6503 12699
rect 15577 12665 15611 12699
rect 18981 12665 19015 12699
rect 1501 12597 1535 12631
rect 3801 12597 3835 12631
rect 4905 12597 4939 12631
rect 6009 12597 6043 12631
rect 6653 12597 6687 12631
rect 7113 12597 7147 12631
rect 11161 12597 11195 12631
rect 14381 12597 14415 12631
rect 18613 12597 18647 12631
rect 21189 12597 21223 12631
rect 24777 12597 24811 12631
rect 6377 12393 6411 12427
rect 7481 12393 7515 12427
rect 11345 12393 11379 12427
rect 14473 12393 14507 12427
rect 18889 12393 18923 12427
rect 19901 12393 19935 12427
rect 23397 12393 23431 12427
rect 25237 12393 25271 12427
rect 10149 12325 10183 12359
rect 1685 12257 1719 12291
rect 4169 12257 4203 12291
rect 4445 12257 4479 12291
rect 10701 12257 10735 12291
rect 11897 12257 11931 12291
rect 13921 12257 13955 12291
rect 14933 12257 14967 12291
rect 15025 12257 15059 12291
rect 16681 12257 16715 12291
rect 20453 12257 20487 12291
rect 23857 12257 23891 12291
rect 1501 12189 1535 12223
rect 2145 12189 2179 12223
rect 2789 12189 2823 12223
rect 4721 12189 4755 12223
rect 5733 12189 5767 12223
rect 6837 12189 6871 12223
rect 7941 12189 7975 12223
rect 9505 12189 9539 12223
rect 11713 12189 11747 12223
rect 14105 12189 14139 12223
rect 14841 12189 14875 12223
rect 16037 12189 16071 12223
rect 17141 12189 17175 12223
rect 18245 12189 18279 12223
rect 20085 12189 20119 12223
rect 22753 12189 22787 12223
rect 24593 12189 24627 12223
rect 3249 12121 3283 12155
rect 9689 12121 9723 12155
rect 10609 12121 10643 12155
rect 12541 12121 12575 12155
rect 13369 12121 13403 12155
rect 20729 12121 20763 12155
rect 1961 12053 1995 12087
rect 2605 12053 2639 12087
rect 3985 12053 4019 12087
rect 8585 12053 8619 12087
rect 9045 12053 9079 12087
rect 10517 12053 10551 12087
rect 11805 12053 11839 12087
rect 15485 12053 15519 12087
rect 15761 12053 15795 12087
rect 17785 12053 17819 12087
rect 19349 12053 19383 12087
rect 19441 12053 19475 12087
rect 19717 12053 19751 12087
rect 22201 12053 22235 12087
rect 1869 11849 1903 11883
rect 2513 11849 2547 11883
rect 5089 11849 5123 11883
rect 9781 11849 9815 11883
rect 10149 11849 10183 11883
rect 10977 11849 11011 11883
rect 11529 11849 11563 11883
rect 11805 11849 11839 11883
rect 12081 11849 12115 11883
rect 13277 11849 13311 11883
rect 13645 11849 13679 11883
rect 13737 11849 13771 11883
rect 14473 11849 14507 11883
rect 14933 11849 14967 11883
rect 16865 11849 16899 11883
rect 17325 11849 17359 11883
rect 21373 11849 21407 11883
rect 4353 11781 4387 11815
rect 4445 11781 4479 11815
rect 6745 11781 6779 11815
rect 10241 11781 10275 11815
rect 18061 11781 18095 11815
rect 19257 11781 19291 11815
rect 23305 11781 23339 11815
rect 1593 11713 1627 11747
rect 2053 11713 2087 11747
rect 2697 11713 2731 11747
rect 3341 11713 3375 11747
rect 3985 11713 4019 11747
rect 5365 11713 5399 11747
rect 12449 11713 12483 11747
rect 12541 11713 12575 11747
rect 14841 11713 14875 11747
rect 15669 11713 15703 11747
rect 17233 11713 17267 11747
rect 19625 11713 19659 11747
rect 20729 11713 20763 11747
rect 22109 11713 22143 11747
rect 23949 11713 23983 11747
rect 6009 11645 6043 11679
rect 7389 11645 7423 11679
rect 7665 11645 7699 11679
rect 10425 11645 10459 11679
rect 12725 11645 12759 11679
rect 13829 11645 13863 11679
rect 15117 11645 15151 11679
rect 17509 11645 17543 11679
rect 18889 11645 18923 11679
rect 24777 11645 24811 11679
rect 6929 11577 6963 11611
rect 9137 11577 9171 11611
rect 3157 11509 3191 11543
rect 3801 11509 3835 11543
rect 9505 11509 9539 11543
rect 16313 11509 16347 11543
rect 20269 11509 20303 11543
rect 1593 11305 1627 11339
rect 4077 11305 4111 11339
rect 7481 11305 7515 11339
rect 8585 11305 8619 11339
rect 10241 11305 10275 11339
rect 11437 11305 11471 11339
rect 13645 11305 13679 11339
rect 13921 11305 13955 11339
rect 14933 11305 14967 11339
rect 17877 11305 17911 11339
rect 18061 11305 18095 11339
rect 19349 11305 19383 11339
rect 19625 11305 19659 11339
rect 25237 11305 25271 11339
rect 2605 11237 2639 11271
rect 22201 11237 22235 11271
rect 2329 11169 2363 11203
rect 5457 11169 5491 11203
rect 10885 11169 10919 11203
rect 11989 11169 12023 11203
rect 13277 11169 13311 11203
rect 15393 11169 15427 11203
rect 16589 11169 16623 11203
rect 17601 11169 17635 11203
rect 18705 11169 18739 11203
rect 19441 11169 19475 11203
rect 20177 11169 20211 11203
rect 1777 11101 1811 11135
rect 2789 11101 2823 11135
rect 4261 11101 4295 11135
rect 4905 11101 4939 11135
rect 5733 11101 5767 11135
rect 6837 11101 6871 11135
rect 7941 11101 7975 11135
rect 9137 11101 9171 11135
rect 10701 11101 10735 11135
rect 11897 11101 11931 11135
rect 14289 11101 14323 11135
rect 16405 11101 16439 11135
rect 16497 11101 16531 11135
rect 17417 11101 17451 11135
rect 20821 11101 20855 11135
rect 22753 11101 22787 11135
rect 24593 11101 24627 11135
rect 2145 11033 2179 11067
rect 3157 11033 3191 11067
rect 3249 11033 3283 11067
rect 5181 11033 5215 11067
rect 9781 11033 9815 11067
rect 13001 11033 13035 11067
rect 13093 11033 13127 11067
rect 18429 11033 18463 11067
rect 21465 11033 21499 11067
rect 22017 11033 22051 11067
rect 23857 11033 23891 11067
rect 4721 10965 4755 10999
rect 6377 10965 6411 10999
rect 10609 10965 10643 10999
rect 11805 10965 11839 10999
rect 12633 10965 12667 10999
rect 16037 10965 16071 10999
rect 18521 10965 18555 10999
rect 19993 10965 20027 10999
rect 20085 10965 20119 10999
rect 1777 10761 1811 10795
rect 8861 10761 8895 10795
rect 12725 10761 12759 10795
rect 13185 10761 13219 10795
rect 15945 10761 15979 10795
rect 16681 10761 16715 10795
rect 18153 10761 18187 10795
rect 21189 10761 21223 10795
rect 25237 10761 25271 10795
rect 3433 10693 3467 10727
rect 7297 10693 7331 10727
rect 7481 10693 7515 10727
rect 9597 10693 9631 10727
rect 12081 10693 12115 10727
rect 14289 10693 14323 10727
rect 15209 10693 15243 10727
rect 20269 10693 20303 10727
rect 22385 10693 22419 10727
rect 23305 10693 23339 10727
rect 25053 10693 25087 10727
rect 1593 10625 1627 10659
rect 2881 10625 2915 10659
rect 4905 10625 4939 10659
rect 5365 10625 5399 10659
rect 6745 10609 6779 10643
rect 8217 10625 8251 10659
rect 13093 10625 13127 10659
rect 17049 10625 17083 10659
rect 18521 10625 18555 10659
rect 19625 10625 19659 10659
rect 21097 10625 21131 10659
rect 22109 10625 22143 10659
rect 23029 10625 23063 10659
rect 2053 10557 2087 10591
rect 3617 10557 3651 10591
rect 4077 10557 4111 10591
rect 9321 10557 9355 10591
rect 13277 10557 13311 10591
rect 14381 10557 14415 10591
rect 14565 10557 14599 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 18613 10557 18647 10591
rect 18797 10557 18831 10591
rect 21281 10557 21315 10591
rect 25421 10557 25455 10591
rect 4721 10489 4755 10523
rect 11069 10489 11103 10523
rect 15577 10489 15611 10523
rect 19257 10489 19291 10523
rect 2697 10421 2731 10455
rect 6009 10421 6043 10455
rect 6561 10421 6595 10455
rect 7941 10421 7975 10455
rect 11713 10421 11747 10455
rect 12173 10421 12207 10455
rect 13921 10421 13955 10455
rect 15025 10421 15059 10455
rect 17693 10421 17727 10455
rect 20729 10421 20763 10455
rect 24777 10421 24811 10455
rect 2973 10217 3007 10251
rect 8585 10217 8619 10251
rect 11253 10217 11287 10251
rect 11805 10217 11839 10251
rect 13001 10217 13035 10251
rect 14736 10217 14770 10251
rect 16681 10217 16715 10251
rect 17785 10217 17819 10251
rect 20085 10217 20119 10251
rect 22845 10217 22879 10251
rect 25237 10217 25271 10251
rect 1593 10149 1627 10183
rect 2237 10149 2271 10183
rect 3985 10149 4019 10183
rect 11437 10149 11471 10183
rect 22385 10149 22419 10183
rect 4721 10081 4755 10115
rect 6377 10081 6411 10115
rect 9137 10081 9171 10115
rect 10885 10081 10919 10115
rect 12357 10081 12391 10115
rect 13553 10081 13587 10115
rect 23489 10081 23523 10115
rect 1777 10013 1811 10047
rect 2421 10013 2455 10047
rect 4169 10013 4203 10047
rect 5733 10013 5767 10047
rect 6837 10013 6871 10047
rect 7941 10013 7975 10047
rect 12173 10013 12207 10047
rect 13369 10013 13403 10047
rect 14473 10013 14507 10047
rect 16589 10013 16623 10047
rect 17141 10013 17175 10047
rect 18245 10013 18279 10047
rect 19441 10013 19475 10047
rect 20637 10013 20671 10047
rect 23213 10013 23247 10047
rect 24593 10013 24627 10047
rect 2789 9945 2823 9979
rect 3249 9945 3283 9979
rect 9413 9945 9447 9979
rect 12265 9945 12299 9979
rect 20913 9945 20947 9979
rect 5273 9877 5307 9911
rect 7481 9877 7515 9911
rect 13461 9877 13495 9911
rect 14197 9877 14231 9911
rect 16221 9877 16255 9911
rect 18889 9877 18923 9911
rect 23305 9877 23339 9911
rect 23857 9877 23891 9911
rect 24041 9877 24075 9911
rect 13461 9673 13495 9707
rect 14565 9673 14599 9707
rect 1409 9605 1443 9639
rect 3249 9605 3283 9639
rect 4169 9605 4203 9639
rect 4721 9605 4755 9639
rect 7297 9605 7331 9639
rect 11345 9605 11379 9639
rect 16129 9605 16163 9639
rect 16957 9605 16991 9639
rect 19625 9605 19659 9639
rect 2145 9537 2179 9571
rect 2797 9537 2831 9571
rect 3985 9537 4019 9571
rect 5365 9537 5399 9571
rect 6009 9537 6043 9571
rect 6653 9537 6687 9571
rect 7757 9537 7791 9571
rect 10885 9537 10919 9571
rect 14933 9537 14967 9571
rect 18153 9537 18187 9571
rect 18981 9537 19015 9571
rect 20269 9537 20303 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 1685 9469 1719 9503
rect 8861 9469 8895 9503
rect 9137 9469 9171 9503
rect 11713 9469 11747 9503
rect 11989 9469 12023 9503
rect 13921 9469 13955 9503
rect 15025 9469 15059 9503
rect 15117 9469 15151 9503
rect 18245 9469 18279 9503
rect 18337 9469 18371 9503
rect 21281 9469 21315 9503
rect 23305 9469 23339 9503
rect 24777 9469 24811 9503
rect 1961 9401 1995 9435
rect 15669 9401 15703 9435
rect 16313 9401 16347 9435
rect 17417 9401 17451 9435
rect 2605 9333 2639 9367
rect 4813 9333 4847 9367
rect 8401 9333 8435 9367
rect 10609 9333 10643 9367
rect 11161 9333 11195 9367
rect 17049 9333 17083 9367
rect 17785 9333 17819 9367
rect 2513 9129 2547 9163
rect 9045 9129 9079 9163
rect 11161 9129 11195 9163
rect 11713 9129 11747 9163
rect 12633 9129 12667 9163
rect 14749 9129 14783 9163
rect 15945 9129 15979 9163
rect 19349 9129 19383 9163
rect 21649 9129 21683 9163
rect 25237 9129 25271 9163
rect 1869 9061 1903 9095
rect 7481 8993 7515 9027
rect 14105 8993 14139 9027
rect 14381 8993 14415 9027
rect 15393 8993 15427 9027
rect 16497 8993 16531 9027
rect 17417 8993 17451 9027
rect 19901 8993 19935 9027
rect 22293 8993 22327 9027
rect 2053 8925 2087 8959
rect 2697 8925 2731 8959
rect 3433 8925 3467 8959
rect 4629 8925 4663 8959
rect 5273 8925 5307 8959
rect 5733 8925 5767 8959
rect 6837 8925 6871 8959
rect 7941 8925 7975 8959
rect 9413 8925 9447 8959
rect 10517 8925 10551 8959
rect 11989 8925 12023 8959
rect 13093 8925 13127 8959
rect 17141 8925 17175 8959
rect 24593 8925 24627 8959
rect 3249 8857 3283 8891
rect 16405 8857 16439 8891
rect 20177 8857 20211 8891
rect 22109 8857 22143 8891
rect 22569 8857 22603 8891
rect 1501 8789 1535 8823
rect 3985 8789 4019 8823
rect 6377 8789 6411 8823
rect 8585 8789 8619 8823
rect 10057 8789 10091 8823
rect 11437 8789 11471 8823
rect 13737 8789 13771 8823
rect 15117 8789 15151 8823
rect 15209 8789 15243 8823
rect 16313 8789 16347 8823
rect 18889 8789 18923 8823
rect 19441 8789 19475 8823
rect 21925 8789 21959 8823
rect 24041 8789 24075 8823
rect 1777 8585 1811 8619
rect 3341 8585 3375 8619
rect 7205 8585 7239 8619
rect 8309 8585 8343 8619
rect 10977 8585 11011 8619
rect 12449 8585 12483 8619
rect 14013 8585 14047 8619
rect 14381 8585 14415 8619
rect 17233 8585 17267 8619
rect 1501 8517 1535 8551
rect 3249 8517 3283 8551
rect 3985 8517 4019 8551
rect 4721 8517 4755 8551
rect 4905 8517 4939 8551
rect 9045 8517 9079 8551
rect 14473 8517 14507 8551
rect 19441 8517 19475 8551
rect 25145 8517 25179 8551
rect 1961 8449 1995 8483
rect 2513 8449 2547 8483
rect 5365 8449 5399 8483
rect 6561 8449 6595 8483
rect 7665 8449 7699 8483
rect 11161 8449 11195 8483
rect 11805 8449 11839 8483
rect 12909 8449 12943 8483
rect 15945 8449 15979 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 20085 8449 20119 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 4169 8381 4203 8415
rect 8769 8381 8803 8415
rect 13921 8381 13955 8415
rect 14565 8381 14599 8415
rect 15209 8381 15243 8415
rect 16037 8381 16071 8415
rect 16221 8381 16255 8415
rect 17325 8381 17359 8415
rect 17417 8381 17451 8415
rect 21281 8381 21315 8415
rect 23305 8381 23339 8415
rect 2697 8313 2731 8347
rect 10517 8313 10551 8347
rect 13553 8313 13587 8347
rect 15025 8313 15059 8347
rect 15577 8313 15611 8347
rect 16865 8313 16899 8347
rect 6009 8245 6043 8279
rect 4813 8041 4847 8075
rect 5273 8041 5307 8075
rect 5457 8041 5491 8075
rect 6377 8041 6411 8075
rect 7481 8041 7515 8075
rect 10701 8041 10735 8075
rect 11161 8041 11195 8075
rect 20453 8041 20487 8075
rect 25237 8041 25271 8075
rect 3433 7973 3467 8007
rect 15669 7973 15703 8007
rect 16865 7973 16899 8007
rect 19441 7973 19475 8007
rect 1501 7905 1535 7939
rect 11621 7905 11655 7939
rect 11805 7905 11839 7939
rect 12909 7905 12943 7939
rect 14841 7905 14875 7939
rect 15393 7905 15427 7939
rect 16221 7905 16255 7939
rect 20085 7905 20119 7939
rect 23857 7905 23891 7939
rect 2513 7837 2547 7871
rect 3249 7837 3283 7871
rect 4721 7837 4755 7871
rect 5733 7837 5767 7871
rect 6837 7837 6871 7871
rect 7941 7837 7975 7871
rect 9045 7837 9079 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 10057 7837 10091 7871
rect 13737 7837 13771 7871
rect 16037 7837 16071 7871
rect 17049 7837 17083 7871
rect 17509 7837 17543 7871
rect 20821 7837 20855 7871
rect 22661 7837 22695 7871
rect 24593 7837 24627 7871
rect 2697 7769 2731 7803
rect 11529 7769 11563 7803
rect 14749 7769 14783 7803
rect 16129 7769 16163 7803
rect 18705 7769 18739 7803
rect 19809 7769 19843 7803
rect 22017 7769 22051 7803
rect 1777 7701 1811 7735
rect 3985 7701 4019 7735
rect 8585 7701 8619 7735
rect 12357 7701 12391 7735
rect 12725 7701 12759 7735
rect 12817 7701 12851 7735
rect 13553 7701 13587 7735
rect 14289 7701 14323 7735
rect 14657 7701 14691 7735
rect 19257 7701 19291 7735
rect 19901 7701 19935 7735
rect 24409 7701 24443 7735
rect 2329 7497 2363 7531
rect 6009 7497 6043 7531
rect 24041 7497 24075 7531
rect 3709 7429 3743 7463
rect 8677 7429 8711 7463
rect 16313 7429 16347 7463
rect 17325 7429 17359 7463
rect 17509 7429 17543 7463
rect 18153 7429 18187 7463
rect 24225 7429 24259 7463
rect 1685 7361 1719 7395
rect 2789 7361 2823 7395
rect 4261 7361 4295 7395
rect 5365 7361 5399 7395
rect 6929 7361 6963 7395
rect 8033 7361 8067 7395
rect 11253 7361 11287 7395
rect 11621 7361 11655 7395
rect 11805 7361 11839 7395
rect 11989 7361 12023 7395
rect 12633 7361 12667 7395
rect 15669 7361 15703 7395
rect 17049 7361 17083 7395
rect 20085 7361 20119 7395
rect 22017 7361 22051 7395
rect 24409 7361 24443 7395
rect 9137 7293 9171 7327
rect 9413 7293 9447 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 13461 7293 13495 7327
rect 13737 7293 13771 7327
rect 17877 7293 17911 7327
rect 21281 7293 21315 7327
rect 24685 7293 24719 7327
rect 3985 7225 4019 7259
rect 10885 7225 10919 7259
rect 23765 7225 23799 7259
rect 3433 7157 3467 7191
rect 4905 7157 4939 7191
rect 6377 7157 6411 7191
rect 6653 7157 6687 7191
rect 7573 7157 7607 7191
rect 12265 7157 12299 7191
rect 15209 7157 15243 7191
rect 16865 7157 16899 7191
rect 19625 7157 19659 7191
rect 22274 7157 22308 7191
rect 8953 6953 8987 6987
rect 1593 6817 1627 6851
rect 9229 6817 9263 6851
rect 10609 6817 10643 6851
rect 12357 6817 12391 6851
rect 12725 6817 12759 6851
rect 15669 6817 15703 6851
rect 18613 6817 18647 6851
rect 19993 6817 20027 6851
rect 20453 6817 20487 6851
rect 25329 6817 25363 6851
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 2881 6749 2915 6783
rect 3985 6749 4019 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 6837 6749 6871 6783
rect 7941 6749 7975 6783
rect 9505 6749 9539 6783
rect 10149 6749 10183 6783
rect 13093 6749 13127 6783
rect 16405 6749 16439 6783
rect 17509 6749 17543 6783
rect 19809 6749 19843 6783
rect 20821 6749 20855 6783
rect 22661 6749 22695 6783
rect 24685 6749 24719 6783
rect 2145 6681 2179 6715
rect 8585 6681 8619 6715
rect 10885 6681 10919 6715
rect 14381 6681 14415 6715
rect 14565 6681 14599 6715
rect 16773 6681 16807 6715
rect 21925 6681 21959 6715
rect 23857 6681 23891 6715
rect 4629 6613 4663 6647
rect 5089 6613 5123 6647
rect 6377 6613 6411 6647
rect 7481 6613 7515 6647
rect 13737 6613 13771 6647
rect 15025 6613 15059 6647
rect 15393 6613 15427 6647
rect 15485 6613 15519 6647
rect 19441 6613 19475 6647
rect 19901 6613 19935 6647
rect 3387 6409 3421 6443
rect 11161 6409 11195 6443
rect 12817 6409 12851 6443
rect 16037 6409 16071 6443
rect 17325 6409 17359 6443
rect 21557 6409 21591 6443
rect 4721 6341 4755 6375
rect 7849 6341 7883 6375
rect 9689 6341 9723 6375
rect 13093 6341 13127 6375
rect 13645 6341 13679 6375
rect 15485 6341 15519 6375
rect 15945 6341 15979 6375
rect 1593 6273 1627 6307
rect 5365 6273 5399 6307
rect 7205 6273 7239 6307
rect 8309 6273 8343 6307
rect 12081 6273 12115 6307
rect 13737 6273 13771 6307
rect 14473 6273 14507 6307
rect 17233 6273 17267 6307
rect 18245 6273 18279 6307
rect 20821 6273 20855 6307
rect 22109 6273 22143 6307
rect 23949 6273 23983 6307
rect 1869 6205 1903 6239
rect 2145 6205 2179 6239
rect 3157 6205 3191 6239
rect 4353 6205 4387 6239
rect 6561 6205 6595 6239
rect 9413 6205 9447 6239
rect 12173 6205 12207 6239
rect 12357 6205 12391 6239
rect 13921 6205 13955 6239
rect 16129 6205 16163 6239
rect 17417 6205 17451 6239
rect 18521 6205 18555 6239
rect 20913 6205 20947 6239
rect 21005 6205 21039 6239
rect 22477 6205 22511 6239
rect 24777 6205 24811 6239
rect 6009 6137 6043 6171
rect 12909 6137 12943 6171
rect 13277 6137 13311 6171
rect 4813 6069 4847 6103
rect 6469 6069 6503 6103
rect 8953 6069 8987 6103
rect 11713 6069 11747 6103
rect 15117 6069 15151 6103
rect 15577 6069 15611 6103
rect 16865 6069 16899 6103
rect 17969 6069 18003 6103
rect 19993 6069 20027 6103
rect 20269 6069 20303 6103
rect 20453 6069 20487 6103
rect 1593 5865 1627 5899
rect 4629 5865 4663 5899
rect 8585 5865 8619 5899
rect 9137 5865 9171 5899
rect 10057 5865 10091 5899
rect 12357 5865 12391 5899
rect 12725 5865 12759 5899
rect 18889 5865 18923 5899
rect 7481 5797 7515 5831
rect 10517 5797 10551 5831
rect 14289 5797 14323 5831
rect 2881 5729 2915 5763
rect 11069 5729 11103 5763
rect 19901 5729 19935 5763
rect 21741 5729 21775 5763
rect 23489 5729 23523 5763
rect 25053 5729 25087 5763
rect 25237 5729 25271 5763
rect 1961 5661 1995 5695
rect 2513 5661 2547 5695
rect 2605 5661 2639 5695
rect 3985 5661 4019 5695
rect 4997 5661 5031 5695
rect 5089 5661 5123 5695
rect 5733 5661 5767 5695
rect 6837 5661 6871 5695
rect 7941 5661 7975 5695
rect 9413 5661 9447 5695
rect 11713 5661 11747 5695
rect 13093 5661 13127 5695
rect 14749 5661 14783 5695
rect 16037 5661 16071 5695
rect 18245 5661 18279 5695
rect 19625 5661 19659 5695
rect 21281 5661 21315 5695
rect 23213 5661 23247 5695
rect 2145 5593 2179 5627
rect 16313 5593 16347 5627
rect 24409 5593 24443 5627
rect 24961 5593 24995 5627
rect 6377 5525 6411 5559
rect 10885 5525 10919 5559
rect 10977 5525 11011 5559
rect 13737 5525 13771 5559
rect 14473 5525 14507 5559
rect 14979 5525 15013 5559
rect 17785 5525 17819 5559
rect 24593 5525 24627 5559
rect 2237 5321 2271 5355
rect 5089 5321 5123 5355
rect 7849 5321 7883 5355
rect 11161 5321 11195 5355
rect 15209 5321 15243 5355
rect 15945 5321 15979 5355
rect 16865 5321 16899 5355
rect 17141 5321 17175 5355
rect 21189 5321 21223 5355
rect 13369 5253 13403 5287
rect 1593 5185 1627 5219
rect 2697 5185 2731 5219
rect 4169 5185 4203 5219
rect 5365 5185 5399 5219
rect 7205 5185 7239 5219
rect 8309 5185 8343 5219
rect 9413 5185 9447 5219
rect 10057 5185 10091 5219
rect 10517 5185 10551 5219
rect 11621 5185 11655 5219
rect 11989 5185 12023 5219
rect 15853 5185 15887 5219
rect 17417 5185 17451 5219
rect 19257 5185 19291 5219
rect 21373 5185 21407 5219
rect 22017 5185 22051 5219
rect 23949 5185 23983 5219
rect 3341 5117 3375 5151
rect 3893 5117 3927 5151
rect 6561 5117 6595 5151
rect 13093 5117 13127 5151
rect 16037 5117 16071 5151
rect 16681 5117 16715 5151
rect 18337 5117 18371 5151
rect 19717 5117 19751 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 6009 4981 6043 5015
rect 8953 4981 8987 5015
rect 12633 4981 12667 5015
rect 14841 4981 14875 5015
rect 15301 4981 15335 5015
rect 15485 4981 15519 5015
rect 7665 4777 7699 4811
rect 8585 4777 8619 4811
rect 9137 4777 9171 4811
rect 22201 4777 22235 4811
rect 14657 4709 14691 4743
rect 19073 4709 19107 4743
rect 1869 4641 1903 4675
rect 5089 4641 5123 4675
rect 15117 4641 15151 4675
rect 16865 4641 16899 4675
rect 20269 4641 20303 4675
rect 20453 4641 20487 4675
rect 23121 4641 23155 4675
rect 1593 4573 1627 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 7113 4573 7147 4607
rect 7941 4573 7975 4607
rect 9321 4573 9355 4607
rect 9781 4573 9815 4607
rect 10885 4573 10919 4607
rect 11989 4573 12023 4607
rect 13093 4573 13127 4607
rect 13737 4573 13771 4607
rect 17325 4573 17359 4607
rect 19441 4573 19475 4607
rect 22661 4573 22695 4607
rect 24593 4573 24627 4607
rect 5365 4505 5399 4539
rect 10425 4505 10459 4539
rect 12633 4505 12667 4539
rect 14473 4505 14507 4539
rect 15393 4505 15427 4539
rect 18429 4505 18463 4539
rect 19717 4505 19751 4539
rect 20729 4505 20763 4539
rect 2881 4437 2915 4471
rect 3341 4437 3375 4471
rect 4629 4437 4663 4471
rect 7481 4437 7515 4471
rect 11529 4437 11563 4471
rect 25237 4437 25271 4471
rect 2881 4233 2915 4267
rect 5457 4233 5491 4267
rect 6561 4233 6595 4267
rect 17417 4233 17451 4267
rect 1593 4097 1627 4131
rect 2789 4097 2823 4131
rect 3065 4097 3099 4131
rect 4813 4097 4847 4131
rect 5825 4097 5859 4131
rect 6745 4097 6779 4131
rect 7205 4097 7239 4131
rect 8309 4097 8343 4131
rect 9413 4097 9447 4131
rect 10517 4097 10551 4131
rect 11529 4097 11563 4131
rect 12173 4097 12207 4131
rect 13369 4097 13403 4131
rect 14013 4097 14047 4131
rect 16221 4097 16255 4131
rect 16405 4097 16439 4131
rect 16773 4097 16807 4131
rect 17509 4097 17543 4131
rect 22201 4097 22235 4131
rect 23857 4097 23891 4131
rect 1869 4029 1903 4063
rect 3525 4029 3559 4063
rect 3801 4029 3835 4063
rect 14289 4029 14323 4063
rect 17601 4029 17635 4063
rect 18245 4029 18279 4063
rect 18521 4029 18555 4063
rect 20361 4029 20395 4063
rect 20637 4029 20671 4063
rect 20913 4029 20947 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 11161 3961 11195 3995
rect 5917 3893 5951 3927
rect 6193 3893 6227 3927
rect 7849 3893 7883 3927
rect 8953 3893 8987 3927
rect 10057 3893 10091 3927
rect 11897 3893 11931 3927
rect 15761 3893 15795 3927
rect 16037 3893 16071 3927
rect 17049 3893 17083 3927
rect 19993 3893 20027 3927
rect 2053 3689 2087 3723
rect 3801 3689 3835 3723
rect 9137 3689 9171 3723
rect 11529 3689 11563 3723
rect 24225 3689 24259 3723
rect 6377 3621 6411 3655
rect 23305 3621 23339 3655
rect 23673 3621 23707 3655
rect 2605 3553 2639 3587
rect 3985 3553 4019 3587
rect 12817 3553 12851 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 18061 3553 18095 3587
rect 19441 3553 19475 3587
rect 22109 3553 22143 3587
rect 23489 3553 23523 3587
rect 1961 3485 1995 3519
rect 2881 3485 2915 3519
rect 4261 3485 4295 3519
rect 5273 3485 5307 3519
rect 6837 3485 6871 3519
rect 7941 3485 7975 3519
rect 9321 3485 9355 3519
rect 9781 3485 9815 3519
rect 10885 3485 10919 3519
rect 12541 3485 12575 3519
rect 14473 3485 14507 3519
rect 16221 3485 16255 3519
rect 18337 3485 18371 3519
rect 21649 3485 21683 3519
rect 24685 3485 24719 3519
rect 1593 3417 1627 3451
rect 6561 3417 6595 3451
rect 11897 3417 11931 3451
rect 19717 3417 19751 3451
rect 25053 3417 25087 3451
rect 5917 3349 5951 3383
rect 7481 3349 7515 3383
rect 8585 3349 8619 3383
rect 10425 3349 10459 3383
rect 11989 3349 12023 3383
rect 21189 3349 21223 3383
rect 23857 3349 23891 3383
rect 6193 3145 6227 3179
rect 6561 3145 6595 3179
rect 8953 3145 8987 3179
rect 10057 3145 10091 3179
rect 1685 3077 1719 3111
rect 1869 3077 1903 3111
rect 11161 3077 11195 3111
rect 2605 3009 2639 3043
rect 3893 3009 3927 3043
rect 4905 3009 4939 3043
rect 5181 3009 5215 3043
rect 6745 3009 6779 3043
rect 7205 3009 7239 3043
rect 8309 3009 8343 3043
rect 9413 3009 9447 3043
rect 10517 3009 10551 3043
rect 13185 3009 13219 3043
rect 15025 3009 15059 3043
rect 16865 3009 16899 3043
rect 18889 3009 18923 3043
rect 20637 3009 20671 3043
rect 20913 3009 20947 3043
rect 22109 3009 22143 3043
rect 23857 3009 23891 3043
rect 2329 2941 2363 2975
rect 3617 2941 3651 2975
rect 6377 2941 6411 2975
rect 7849 2941 7883 2975
rect 11713 2941 11747 2975
rect 11989 2941 12023 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 22477 2941 22511 2975
rect 24317 2941 24351 2975
rect 3525 2873 3559 2907
rect 1501 2601 1535 2635
rect 2053 2601 2087 2635
rect 9137 2601 9171 2635
rect 23765 2601 23799 2635
rect 24041 2601 24075 2635
rect 25237 2601 25271 2635
rect 4629 2533 4663 2567
rect 7205 2533 7239 2567
rect 24225 2533 24259 2567
rect 2605 2465 2639 2499
rect 5457 2465 5491 2499
rect 11713 2465 11747 2499
rect 14933 2465 14967 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 1961 2397 1995 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 5181 2397 5215 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 8033 2397 8067 2431
rect 9321 2397 9355 2431
rect 9781 2397 9815 2431
rect 12541 2397 12575 2431
rect 14657 2397 14691 2431
rect 17049 2397 17083 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 21465 2397 21499 2431
rect 22017 2397 22051 2431
rect 24593 2397 24627 2431
rect 10977 2329 11011 2363
rect 13277 2329 13311 2363
rect 16405 2329 16439 2363
rect 7665 2261 7699 2295
rect 14105 2261 14139 2295
rect 16129 2261 16163 2295
rect 18705 2261 18739 2295
rect 21097 2261 21131 2295
rect 21281 2261 21315 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 18966 54272 18972 54324
rect 19024 54272 19030 54324
rect 18141 54247 18199 54253
rect 18141 54244 18153 54247
rect 17880 54216 18153 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 3878 54176 3884 54188
rect 2271 54148 3884 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 3878 54136 3884 54148
rect 3936 54136 3942 54188
rect 4157 54179 4215 54185
rect 4157 54145 4169 54179
rect 4203 54176 4215 54179
rect 6546 54176 6552 54188
rect 4203 54148 6552 54176
rect 4203 54145 4215 54148
rect 4157 54139 4215 54145
rect 6546 54136 6552 54148
rect 6604 54136 6610 54188
rect 6730 54136 6736 54188
rect 6788 54136 6794 54188
rect 13446 54136 13452 54188
rect 13504 54176 13510 54188
rect 13725 54179 13783 54185
rect 13725 54176 13737 54179
rect 13504 54148 13737 54176
rect 13504 54136 13510 54148
rect 13725 54145 13737 54148
rect 13771 54176 13783 54179
rect 14093 54179 14151 54185
rect 14093 54176 14105 54179
rect 13771 54148 14105 54176
rect 13771 54145 13783 54148
rect 13725 54139 13783 54145
rect 14093 54145 14105 54148
rect 14139 54145 14151 54179
rect 14093 54139 14151 54145
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15105 54179 15163 54185
rect 15105 54176 15117 54179
rect 14884 54148 15117 54176
rect 14884 54136 14890 54148
rect 15105 54145 15117 54148
rect 15151 54176 15163 54179
rect 15381 54179 15439 54185
rect 15381 54176 15393 54179
rect 15151 54148 15393 54176
rect 15151 54145 15163 54148
rect 15105 54139 15163 54145
rect 15381 54145 15393 54148
rect 15427 54145 15439 54179
rect 15381 54139 15439 54145
rect 16574 54136 16580 54188
rect 16632 54176 16638 54188
rect 17037 54179 17095 54185
rect 17037 54176 17049 54179
rect 16632 54148 17049 54176
rect 16632 54136 16638 54148
rect 17037 54145 17049 54148
rect 17083 54176 17095 54179
rect 17313 54179 17371 54185
rect 17313 54176 17325 54179
rect 17083 54148 17325 54176
rect 17083 54145 17095 54148
rect 17037 54139 17095 54145
rect 17313 54145 17325 54148
rect 17359 54145 17371 54179
rect 17313 54139 17371 54145
rect 17586 54136 17592 54188
rect 17644 54176 17650 54188
rect 17880 54185 17908 54216
rect 18141 54213 18153 54216
rect 18187 54213 18199 54247
rect 25314 54244 25320 54256
rect 18141 54207 18199 54213
rect 22296 54216 25320 54244
rect 22296 54185 22324 54216
rect 25314 54204 25320 54216
rect 25372 54204 25378 54256
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17644 54148 17877 54176
rect 17644 54136 17650 54148
rect 17865 54145 17877 54148
rect 17911 54145 17923 54179
rect 19705 54179 19763 54185
rect 19705 54176 19717 54179
rect 17865 54139 17923 54145
rect 18156 54148 19717 54176
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 4062 54068 4068 54120
rect 4120 54108 4126 54120
rect 4433 54111 4491 54117
rect 4433 54108 4445 54111
rect 4120 54080 4445 54108
rect 4120 54068 4126 54080
rect 4433 54077 4445 54080
rect 4479 54077 4491 54111
rect 4433 54071 4491 54077
rect 6914 54068 6920 54120
rect 6972 54108 6978 54120
rect 7101 54111 7159 54117
rect 7101 54108 7113 54111
rect 6972 54080 7113 54108
rect 6972 54068 6978 54080
rect 7101 54077 7113 54080
rect 7147 54077 7159 54111
rect 7101 54071 7159 54077
rect 11054 54068 11060 54120
rect 11112 54108 11118 54120
rect 18156 54108 18184 54148
rect 19705 54145 19717 54148
rect 19751 54145 19763 54179
rect 19705 54139 19763 54145
rect 21177 54179 21235 54185
rect 21177 54145 21189 54179
rect 21223 54176 21235 54179
rect 22281 54179 22339 54185
rect 21223 54148 21956 54176
rect 21223 54145 21235 54148
rect 21177 54139 21235 54145
rect 11112 54080 18184 54108
rect 11112 54068 11118 54080
rect 18966 54068 18972 54120
rect 19024 54108 19030 54120
rect 19429 54111 19487 54117
rect 19429 54108 19441 54111
rect 19024 54080 19441 54108
rect 19024 54068 19030 54080
rect 19429 54077 19441 54080
rect 19475 54077 19487 54111
rect 19429 54071 19487 54077
rect 16758 54000 16764 54052
rect 16816 54040 16822 54052
rect 21928 54049 21956 54148
rect 22281 54145 22293 54179
rect 22327 54145 22339 54179
rect 22281 54139 22339 54145
rect 23385 54179 23443 54185
rect 23385 54145 23397 54179
rect 23431 54145 23443 54179
rect 23385 54139 23443 54145
rect 24581 54179 24639 54185
rect 24581 54145 24593 54179
rect 24627 54176 24639 54179
rect 25222 54176 25228 54188
rect 24627 54148 25228 54176
rect 24627 54145 24639 54148
rect 24581 54139 24639 54145
rect 23400 54108 23428 54139
rect 25222 54136 25228 54148
rect 25280 54136 25286 54188
rect 25130 54108 25136 54120
rect 23400 54080 25136 54108
rect 25130 54068 25136 54080
rect 25188 54068 25194 54120
rect 21361 54043 21419 54049
rect 21361 54040 21373 54043
rect 16816 54012 21373 54040
rect 16816 54000 16822 54012
rect 21361 54009 21373 54012
rect 21407 54009 21419 54043
rect 21361 54003 21419 54009
rect 21913 54043 21971 54049
rect 21913 54009 21925 54043
rect 21959 54040 21971 54043
rect 23382 54040 23388 54052
rect 21959 54012 23388 54040
rect 21959 54009 21971 54012
rect 21913 54003 21971 54009
rect 23382 54000 23388 54012
rect 23440 54000 23446 54052
rect 23474 54000 23480 54052
rect 23532 54040 23538 54052
rect 25225 54043 25283 54049
rect 25225 54040 25237 54043
rect 23532 54012 25237 54040
rect 23532 54000 23538 54012
rect 25225 54009 25237 54012
rect 25271 54009 25283 54043
rect 25225 54003 25283 54009
rect 13538 53932 13544 53984
rect 13596 53932 13602 53984
rect 14918 53932 14924 53984
rect 14976 53932 14982 53984
rect 15654 53932 15660 53984
rect 15712 53972 15718 53984
rect 16853 53975 16911 53981
rect 16853 53972 16865 53975
rect 15712 53944 16865 53972
rect 15712 53932 15718 53944
rect 16853 53941 16865 53944
rect 16899 53941 16911 53975
rect 16853 53935 16911 53941
rect 17126 53932 17132 53984
rect 17184 53972 17190 53984
rect 17681 53975 17739 53981
rect 17681 53972 17693 53975
rect 17184 53944 17693 53972
rect 17184 53932 17190 53944
rect 17681 53941 17693 53944
rect 17727 53941 17739 53975
rect 17681 53935 17739 53941
rect 22925 53975 22983 53981
rect 22925 53941 22937 53975
rect 22971 53972 22983 53975
rect 23934 53972 23940 53984
rect 22971 53944 23940 53972
rect 22971 53941 22983 53944
rect 22925 53935 22983 53941
rect 23934 53932 23940 53944
rect 23992 53932 23998 53984
rect 24029 53975 24087 53981
rect 24029 53941 24041 53975
rect 24075 53972 24087 53975
rect 24578 53972 24584 53984
rect 24075 53944 24584 53972
rect 24075 53941 24087 53944
rect 24029 53935 24087 53941
rect 24578 53932 24584 53944
rect 24636 53932 24642 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 25222 53728 25228 53780
rect 25280 53728 25286 53780
rect 24213 53703 24271 53709
rect 24213 53669 24225 53703
rect 24259 53700 24271 53703
rect 24854 53700 24860 53712
rect 24259 53672 24860 53700
rect 24259 53669 24271 53672
rect 24213 53663 24271 53669
rect 24854 53660 24860 53672
rect 24912 53700 24918 53712
rect 25866 53700 25872 53712
rect 24912 53672 25872 53700
rect 24912 53660 24918 53672
rect 25866 53660 25872 53672
rect 25924 53660 25930 53712
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 2041 53635 2099 53641
rect 2041 53632 2053 53635
rect 1084 53604 2053 53632
rect 1084 53592 1090 53604
rect 2041 53601 2053 53604
rect 2087 53601 2099 53635
rect 2041 53595 2099 53601
rect 5166 53592 5172 53644
rect 5224 53632 5230 53644
rect 5721 53635 5779 53641
rect 5721 53632 5733 53635
rect 5224 53604 5733 53632
rect 5224 53592 5230 53604
rect 5721 53601 5733 53604
rect 5767 53601 5779 53635
rect 5721 53595 5779 53601
rect 1765 53567 1823 53573
rect 1765 53533 1777 53567
rect 1811 53533 1823 53567
rect 1765 53527 1823 53533
rect 5445 53567 5503 53573
rect 5445 53533 5457 53567
rect 5491 53564 5503 53567
rect 7650 53564 7656 53576
rect 5491 53536 7656 53564
rect 5491 53533 5503 53536
rect 5445 53527 5503 53533
rect 1780 53496 1808 53527
rect 7650 53524 7656 53536
rect 7708 53524 7714 53576
rect 22097 53567 22155 53573
rect 22097 53533 22109 53567
rect 22143 53564 22155 53567
rect 22370 53564 22376 53576
rect 22143 53536 22376 53564
rect 22143 53533 22155 53536
rect 22097 53527 22155 53533
rect 22370 53524 22376 53536
rect 22428 53524 22434 53576
rect 23109 53567 23167 53573
rect 23109 53533 23121 53567
rect 23155 53564 23167 53567
rect 23290 53564 23296 53576
rect 23155 53536 23296 53564
rect 23155 53533 23167 53536
rect 23109 53527 23167 53533
rect 23290 53524 23296 53536
rect 23348 53524 23354 53576
rect 24578 53524 24584 53576
rect 24636 53524 24642 53576
rect 5534 53496 5540 53508
rect 1780 53468 5540 53496
rect 5534 53456 5540 53468
rect 5592 53456 5598 53508
rect 22094 53388 22100 53440
rect 22152 53428 22158 53440
rect 22557 53431 22615 53437
rect 22557 53428 22569 53431
rect 22152 53400 22569 53428
rect 22152 53388 22158 53400
rect 22557 53397 22569 53400
rect 22603 53397 22615 53431
rect 22557 53391 22615 53397
rect 23750 53388 23756 53440
rect 23808 53388 23814 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 3878 53184 3884 53236
rect 3936 53224 3942 53236
rect 4985 53227 5043 53233
rect 4985 53224 4997 53227
rect 3936 53196 4997 53224
rect 3936 53184 3942 53196
rect 4985 53193 4997 53196
rect 5031 53193 5043 53227
rect 4985 53187 5043 53193
rect 6546 53184 6552 53236
rect 6604 53184 6610 53236
rect 25130 53184 25136 53236
rect 25188 53224 25194 53236
rect 25225 53227 25283 53233
rect 25225 53224 25237 53227
rect 25188 53196 25237 53224
rect 25188 53184 25194 53196
rect 25225 53193 25237 53196
rect 25271 53193 25283 53227
rect 25225 53187 25283 53193
rect 22465 53159 22523 53165
rect 22465 53125 22477 53159
rect 22511 53156 22523 53159
rect 22830 53156 22836 53168
rect 22511 53128 22836 53156
rect 22511 53125 22523 53128
rect 22465 53119 22523 53125
rect 22830 53116 22836 53128
rect 22888 53116 22894 53168
rect 24854 53156 24860 53168
rect 23492 53128 24860 53156
rect 5169 53091 5227 53097
rect 5169 53057 5181 53091
rect 5215 53057 5227 53091
rect 5169 53051 5227 53057
rect 6733 53091 6791 53097
rect 6733 53057 6745 53091
rect 6779 53088 6791 53091
rect 8846 53088 8852 53100
rect 6779 53060 8852 53088
rect 6779 53057 6791 53060
rect 6733 53051 6791 53057
rect 5184 53020 5212 53051
rect 8846 53048 8852 53060
rect 8904 53048 8910 53100
rect 16206 53048 16212 53100
rect 16264 53088 16270 53100
rect 20346 53088 20352 53100
rect 16264 53060 20352 53088
rect 16264 53048 16270 53060
rect 20346 53048 20352 53060
rect 20404 53048 20410 53100
rect 23492 53097 23520 53128
rect 24854 53116 24860 53128
rect 24912 53116 24918 53168
rect 23477 53091 23535 53097
rect 23477 53057 23489 53091
rect 23523 53057 23535 53091
rect 23477 53051 23535 53057
rect 23934 53048 23940 53100
rect 23992 53088 23998 53100
rect 24581 53091 24639 53097
rect 24581 53088 24593 53091
rect 23992 53060 24593 53088
rect 23992 53048 23998 53060
rect 24581 53057 24593 53060
rect 24627 53057 24639 53091
rect 24581 53051 24639 53057
rect 7742 53020 7748 53032
rect 5184 52992 7748 53020
rect 7742 52980 7748 52992
rect 7800 52980 7806 53032
rect 18966 52912 18972 52964
rect 19024 52952 19030 52964
rect 23017 52955 23075 52961
rect 23017 52952 23029 52955
rect 19024 52924 23029 52952
rect 19024 52912 19030 52924
rect 23017 52921 23029 52924
rect 23063 52921 23075 52955
rect 23017 52915 23075 52921
rect 24121 52887 24179 52893
rect 24121 52853 24133 52887
rect 24167 52884 24179 52887
rect 24670 52884 24676 52896
rect 24167 52856 24676 52884
rect 24167 52853 24179 52856
rect 24121 52847 24179 52853
rect 24670 52844 24676 52856
rect 24728 52844 24734 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 7650 52640 7656 52692
rect 7708 52640 7714 52692
rect 23109 52683 23167 52689
rect 23109 52649 23121 52683
rect 23155 52680 23167 52683
rect 23290 52680 23296 52692
rect 23155 52652 23296 52680
rect 23155 52649 23167 52652
rect 23109 52643 23167 52649
rect 23290 52640 23296 52652
rect 23348 52640 23354 52692
rect 25314 52640 25320 52692
rect 25372 52640 25378 52692
rect 7834 52572 7840 52624
rect 7892 52612 7898 52624
rect 8386 52612 8392 52624
rect 7892 52584 8392 52612
rect 7892 52572 7898 52584
rect 8386 52572 8392 52584
rect 8444 52572 8450 52624
rect 7837 52479 7895 52485
rect 7837 52445 7849 52479
rect 7883 52476 7895 52479
rect 9582 52476 9588 52488
rect 7883 52448 9588 52476
rect 7883 52445 7895 52448
rect 7837 52439 7895 52445
rect 9582 52436 9588 52448
rect 9640 52436 9646 52488
rect 17218 52436 17224 52488
rect 17276 52476 17282 52488
rect 22738 52476 22744 52488
rect 17276 52448 22744 52476
rect 17276 52436 17282 52448
rect 22738 52436 22744 52448
rect 22796 52436 22802 52488
rect 23293 52479 23351 52485
rect 23293 52445 23305 52479
rect 23339 52476 23351 52479
rect 23474 52476 23480 52488
rect 23339 52448 23480 52476
rect 23339 52445 23351 52448
rect 23293 52439 23351 52445
rect 23474 52436 23480 52448
rect 23532 52436 23538 52488
rect 23753 52479 23811 52485
rect 23753 52445 23765 52479
rect 23799 52476 23811 52479
rect 24118 52476 24124 52488
rect 23799 52448 24124 52476
rect 23799 52445 23811 52448
rect 23753 52439 23811 52445
rect 24118 52436 24124 52448
rect 24176 52436 24182 52488
rect 24670 52436 24676 52488
rect 24728 52436 24734 52488
rect 23934 52300 23940 52352
rect 23992 52300 23998 52352
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 6730 52096 6736 52148
rect 6788 52136 6794 52148
rect 8849 52139 8907 52145
rect 8849 52136 8861 52139
rect 6788 52108 8861 52136
rect 6788 52096 6794 52108
rect 8849 52105 8861 52108
rect 8895 52105 8907 52139
rect 8849 52099 8907 52105
rect 24946 52028 24952 52080
rect 25004 52028 25010 52080
rect 8757 52003 8815 52009
rect 8757 51969 8769 52003
rect 8803 52000 8815 52003
rect 10778 52000 10784 52012
rect 8803 51972 10784 52000
rect 8803 51969 8815 51972
rect 8757 51963 8815 51969
rect 10778 51960 10784 51972
rect 10836 51960 10842 52012
rect 22925 52003 22983 52009
rect 22925 51969 22937 52003
rect 22971 52000 22983 52003
rect 23750 52000 23756 52012
rect 22971 51972 23756 52000
rect 22971 51969 22983 51972
rect 22925 51963 22983 51969
rect 23750 51960 23756 51972
rect 23808 51960 23814 52012
rect 24121 52003 24179 52009
rect 24121 51969 24133 52003
rect 24167 52000 24179 52003
rect 24578 52000 24584 52012
rect 24167 51972 24584 52000
rect 24167 51969 24179 51972
rect 24121 51963 24179 51969
rect 24578 51960 24584 51972
rect 24636 51960 24642 52012
rect 18690 51892 18696 51944
rect 18748 51932 18754 51944
rect 25225 51935 25283 51941
rect 25225 51932 25237 51935
rect 18748 51904 25237 51932
rect 18748 51892 18754 51904
rect 25225 51901 25237 51904
rect 25271 51901 25283 51935
rect 25225 51895 25283 51901
rect 17310 51824 17316 51876
rect 17368 51864 17374 51876
rect 24305 51867 24363 51873
rect 24305 51864 24317 51867
rect 17368 51836 24317 51864
rect 17368 51824 17374 51836
rect 24305 51833 24317 51836
rect 24351 51833 24363 51867
rect 24305 51827 24363 51833
rect 22554 51756 22560 51808
rect 22612 51796 22618 51808
rect 23569 51799 23627 51805
rect 23569 51796 23581 51799
rect 22612 51768 23581 51796
rect 22612 51756 22618 51768
rect 23569 51765 23581 51768
rect 23615 51765 23627 51799
rect 23569 51759 23627 51765
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 24118 51552 24124 51604
rect 24176 51552 24182 51604
rect 24578 51552 24584 51604
rect 24636 51552 24642 51604
rect 23845 51527 23903 51533
rect 23845 51493 23857 51527
rect 23891 51524 23903 51527
rect 24946 51524 24952 51536
rect 23891 51496 24952 51524
rect 23891 51493 23903 51496
rect 23845 51487 23903 51493
rect 24946 51484 24952 51496
rect 25004 51484 25010 51536
rect 24029 51323 24087 51329
rect 24029 51289 24041 51323
rect 24075 51320 24087 51323
rect 24946 51320 24952 51332
rect 24075 51292 24952 51320
rect 24075 51289 24087 51292
rect 24029 51283 24087 51289
rect 24946 51280 24952 51292
rect 25004 51280 25010 51332
rect 25038 51212 25044 51264
rect 25096 51212 25102 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 7742 51008 7748 51060
rect 7800 51048 7806 51060
rect 7929 51051 7987 51057
rect 7929 51048 7941 51051
rect 7800 51020 7941 51048
rect 7800 51008 7806 51020
rect 7929 51017 7941 51020
rect 7975 51017 7987 51051
rect 7929 51011 7987 51017
rect 7469 50915 7527 50921
rect 7469 50881 7481 50915
rect 7515 50912 7527 50915
rect 24581 50915 24639 50921
rect 7515 50884 8432 50912
rect 7515 50881 7527 50884
rect 7469 50875 7527 50881
rect 5534 50668 5540 50720
rect 5592 50708 5598 50720
rect 6822 50708 6828 50720
rect 5592 50680 6828 50708
rect 5592 50668 5598 50680
rect 6822 50668 6828 50680
rect 6880 50708 6886 50720
rect 8404 50717 8432 50884
rect 24581 50881 24593 50915
rect 24627 50912 24639 50915
rect 24946 50912 24952 50924
rect 24627 50884 24952 50912
rect 24627 50881 24639 50884
rect 24581 50875 24639 50881
rect 24946 50872 24952 50884
rect 25004 50872 25010 50924
rect 7561 50711 7619 50717
rect 7561 50708 7573 50711
rect 6880 50680 7573 50708
rect 6880 50668 6886 50680
rect 7561 50677 7573 50680
rect 7607 50677 7619 50711
rect 7561 50671 7619 50677
rect 8389 50711 8447 50717
rect 8389 50677 8401 50711
rect 8435 50708 8447 50711
rect 11054 50708 11060 50720
rect 8435 50680 11060 50708
rect 8435 50677 8447 50680
rect 8389 50671 8447 50677
rect 11054 50668 11060 50680
rect 11112 50668 11118 50720
rect 24578 50668 24584 50720
rect 24636 50708 24642 50720
rect 25041 50711 25099 50717
rect 25041 50708 25053 50711
rect 24636 50680 25053 50708
rect 24636 50668 24642 50680
rect 25041 50677 25053 50680
rect 25087 50677 25099 50711
rect 25041 50671 25099 50677
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 16390 50464 16396 50516
rect 16448 50504 16454 50516
rect 24578 50504 24584 50516
rect 16448 50476 24584 50504
rect 16448 50464 16454 50476
rect 24578 50464 24584 50476
rect 24636 50464 24642 50516
rect 6822 50328 6828 50380
rect 6880 50368 6886 50380
rect 8294 50368 8300 50380
rect 6880 50340 8300 50368
rect 6880 50328 6886 50340
rect 8294 50328 8300 50340
rect 8352 50328 8358 50380
rect 16482 50328 16488 50380
rect 16540 50368 16546 50380
rect 24486 50368 24492 50380
rect 16540 50340 24492 50368
rect 16540 50328 16546 50340
rect 24486 50328 24492 50340
rect 24544 50328 24550 50380
rect 25498 50124 25504 50176
rect 25556 50124 25562 50176
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 24489 49827 24547 49833
rect 24489 49793 24501 49827
rect 24535 49824 24547 49827
rect 25498 49824 25504 49836
rect 24535 49796 25504 49824
rect 24535 49793 24547 49796
rect 24489 49787 24547 49793
rect 25498 49784 25504 49796
rect 25556 49784 25562 49836
rect 24762 49716 24768 49768
rect 24820 49716 24826 49768
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 18782 49376 18788 49428
rect 18840 49416 18846 49428
rect 22094 49416 22100 49428
rect 18840 49388 22100 49416
rect 18840 49376 18846 49388
rect 22094 49376 22100 49388
rect 22152 49376 22158 49428
rect 22554 49172 22560 49224
rect 22612 49172 22618 49224
rect 24765 49147 24823 49153
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 25130 49144 25136 49156
rect 24811 49116 25136 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 25130 49104 25136 49116
rect 25188 49104 25194 49156
rect 22646 49036 22652 49088
rect 22704 49076 22710 49088
rect 23201 49079 23259 49085
rect 23201 49076 23213 49079
rect 22704 49048 23213 49076
rect 22704 49036 22710 49048
rect 23201 49045 23213 49048
rect 23247 49045 23259 49079
rect 23201 49039 23259 49045
rect 25222 49036 25228 49088
rect 25280 49036 25286 49088
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 8846 48832 8852 48884
rect 8904 48872 8910 48884
rect 10505 48875 10563 48881
rect 10505 48872 10517 48875
rect 8904 48844 10517 48872
rect 8904 48832 8910 48844
rect 10505 48841 10517 48844
rect 10551 48872 10563 48875
rect 11422 48872 11428 48884
rect 10551 48844 11428 48872
rect 10551 48841 10563 48844
rect 10505 48835 10563 48841
rect 11422 48832 11428 48844
rect 11480 48832 11486 48884
rect 7742 48764 7748 48816
rect 7800 48804 7806 48816
rect 7929 48807 7987 48813
rect 7929 48804 7941 48807
rect 7800 48776 7941 48804
rect 7800 48764 7806 48776
rect 7929 48773 7941 48776
rect 7975 48804 7987 48807
rect 8202 48804 8208 48816
rect 7975 48776 8208 48804
rect 7975 48773 7987 48776
rect 7929 48767 7987 48773
rect 8202 48764 8208 48776
rect 8260 48764 8266 48816
rect 10965 48807 11023 48813
rect 10965 48773 10977 48807
rect 11011 48804 11023 48807
rect 11054 48804 11060 48816
rect 11011 48776 11060 48804
rect 11011 48773 11023 48776
rect 10965 48767 11023 48773
rect 10045 48739 10103 48745
rect 10045 48705 10057 48739
rect 10091 48736 10103 48739
rect 10980 48736 11008 48767
rect 11054 48764 11060 48776
rect 11112 48764 11118 48816
rect 10091 48708 11008 48736
rect 10091 48705 10103 48708
rect 10045 48699 10103 48705
rect 7742 48628 7748 48680
rect 7800 48628 7806 48680
rect 8386 48628 8392 48680
rect 8444 48628 8450 48680
rect 10134 48492 10140 48544
rect 10192 48492 10198 48544
rect 25130 48492 25136 48544
rect 25188 48532 25194 48544
rect 25409 48535 25467 48541
rect 25409 48532 25421 48535
rect 25188 48504 25421 48532
rect 25188 48492 25194 48504
rect 25409 48501 25421 48504
rect 25455 48501 25467 48535
rect 25409 48495 25467 48501
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 8294 48220 8300 48272
rect 8352 48220 8358 48272
rect 6549 48195 6607 48201
rect 6549 48161 6561 48195
rect 6595 48192 6607 48195
rect 8570 48192 8576 48204
rect 6595 48164 8576 48192
rect 6595 48161 6607 48164
rect 6549 48155 6607 48161
rect 8570 48152 8576 48164
rect 8628 48152 8634 48204
rect 9048 48164 9260 48192
rect 8202 48084 8208 48136
rect 8260 48124 8266 48136
rect 9048 48124 9076 48164
rect 8260 48096 9076 48124
rect 8260 48084 8266 48096
rect 9122 48084 9128 48136
rect 9180 48084 9186 48136
rect 9232 48124 9260 48164
rect 10264 48127 10322 48133
rect 10264 48124 10276 48127
rect 9232 48096 10276 48124
rect 10264 48093 10276 48096
rect 10310 48093 10322 48127
rect 10264 48087 10322 48093
rect 11422 48084 11428 48136
rect 11480 48133 11486 48136
rect 11480 48127 11518 48133
rect 11506 48093 11518 48127
rect 11480 48087 11518 48093
rect 11480 48084 11486 48087
rect 25130 48084 25136 48136
rect 25188 48084 25194 48136
rect 6825 48059 6883 48065
rect 6825 48025 6837 48059
rect 6871 48025 6883 48059
rect 6825 48019 6883 48025
rect 6840 47988 6868 48019
rect 7834 48016 7840 48068
rect 7892 48016 7898 48068
rect 9769 48059 9827 48065
rect 9769 48056 9781 48059
rect 8220 48028 9781 48056
rect 8220 47988 8248 48028
rect 9769 48025 9781 48028
rect 9815 48025 9827 48059
rect 9769 48019 9827 48025
rect 6840 47960 8248 47988
rect 8570 47948 8576 48000
rect 8628 47948 8634 48000
rect 10367 47991 10425 47997
rect 10367 47957 10379 47991
rect 10413 47988 10425 47991
rect 11422 47988 11428 48000
rect 10413 47960 11428 47988
rect 10413 47957 10425 47960
rect 10367 47951 10425 47957
rect 11422 47948 11428 47960
rect 11480 47948 11486 48000
rect 11563 47991 11621 47997
rect 11563 47957 11575 47991
rect 11609 47988 11621 47991
rect 14458 47988 14464 48000
rect 11609 47960 14464 47988
rect 11609 47957 11621 47960
rect 11563 47951 11621 47957
rect 14458 47948 14464 47960
rect 14516 47948 14522 48000
rect 24854 47948 24860 48000
rect 24912 47988 24918 48000
rect 25225 47991 25283 47997
rect 25225 47988 25237 47991
rect 24912 47960 25237 47988
rect 24912 47948 24918 47960
rect 25225 47957 25237 47960
rect 25271 47957 25283 47991
rect 25225 47951 25283 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 8846 47676 8852 47728
rect 8904 47676 8910 47728
rect 12472 47651 12530 47657
rect 12472 47648 12484 47651
rect 10152 47620 12484 47648
rect 8665 47583 8723 47589
rect 8665 47549 8677 47583
rect 8711 47580 8723 47583
rect 8711 47552 8800 47580
rect 8711 47549 8723 47552
rect 8665 47543 8723 47549
rect 8772 47524 8800 47552
rect 9306 47540 9312 47592
rect 9364 47540 9370 47592
rect 9582 47540 9588 47592
rect 9640 47580 9646 47592
rect 10152 47580 10180 47620
rect 12472 47617 12484 47620
rect 12518 47617 12530 47651
rect 12472 47611 12530 47617
rect 24857 47651 24915 47657
rect 24857 47617 24869 47651
rect 24903 47648 24915 47651
rect 25314 47648 25320 47660
rect 24903 47620 25320 47648
rect 24903 47617 24915 47620
rect 24857 47611 24915 47617
rect 25314 47608 25320 47620
rect 25372 47608 25378 47660
rect 9640 47552 10180 47580
rect 9640 47540 9646 47552
rect 8754 47472 8760 47524
rect 8812 47472 8818 47524
rect 7834 47404 7840 47456
rect 7892 47444 7898 47456
rect 8389 47447 8447 47453
rect 8389 47444 8401 47447
rect 7892 47416 8401 47444
rect 7892 47404 7898 47416
rect 8389 47413 8401 47416
rect 8435 47444 8447 47447
rect 10502 47444 10508 47456
rect 8435 47416 10508 47444
rect 8435 47413 8447 47416
rect 8389 47407 8447 47413
rect 10502 47404 10508 47416
rect 10560 47404 10566 47456
rect 12575 47447 12633 47453
rect 12575 47413 12587 47447
rect 12621 47444 12633 47447
rect 14642 47444 14648 47456
rect 12621 47416 14648 47444
rect 12621 47413 12633 47416
rect 12575 47407 12633 47413
rect 14642 47404 14648 47416
rect 14700 47404 14706 47456
rect 25133 47447 25191 47453
rect 25133 47413 25145 47447
rect 25179 47444 25191 47447
rect 25774 47444 25780 47456
rect 25179 47416 25780 47444
rect 25179 47413 25191 47416
rect 25133 47407 25191 47413
rect 25774 47404 25780 47416
rect 25832 47404 25838 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 9122 47200 9128 47252
rect 9180 47240 9186 47252
rect 9769 47243 9827 47249
rect 9769 47240 9781 47243
rect 9180 47212 9781 47240
rect 9180 47200 9186 47212
rect 9769 47209 9781 47212
rect 9815 47209 9827 47243
rect 9769 47203 9827 47209
rect 10318 47200 10324 47252
rect 10376 47200 10382 47252
rect 11054 47200 11060 47252
rect 11112 47200 11118 47252
rect 9582 47132 9588 47184
rect 9640 47172 9646 47184
rect 10689 47175 10747 47181
rect 10689 47172 10701 47175
rect 9640 47144 10701 47172
rect 9640 47132 9646 47144
rect 10689 47141 10701 47144
rect 10735 47141 10747 47175
rect 10689 47135 10747 47141
rect 14277 47107 14335 47113
rect 14277 47073 14289 47107
rect 14323 47104 14335 47107
rect 14918 47104 14924 47116
rect 14323 47076 14924 47104
rect 14323 47073 14335 47076
rect 14277 47067 14335 47073
rect 14918 47064 14924 47076
rect 14976 47064 14982 47116
rect 9125 47039 9183 47045
rect 9125 47005 9137 47039
rect 9171 47036 9183 47039
rect 9766 47036 9772 47048
rect 9171 47008 9772 47036
rect 9171 47005 9183 47008
rect 9125 46999 9183 47005
rect 9766 46996 9772 47008
rect 9824 46996 9830 47048
rect 10229 47039 10287 47045
rect 10229 47005 10241 47039
rect 10275 47036 10287 47039
rect 11054 47036 11060 47048
rect 10275 47008 11060 47036
rect 10275 47005 10287 47008
rect 10229 46999 10287 47005
rect 11054 46996 11060 47008
rect 11112 46996 11118 47048
rect 12158 46996 12164 47048
rect 12216 47036 12222 47048
rect 13300 47039 13358 47045
rect 13300 47036 13312 47039
rect 12216 47008 13312 47036
rect 12216 46996 12222 47008
rect 13300 47005 13312 47008
rect 13346 47005 13358 47039
rect 13300 46999 13358 47005
rect 22646 46996 22652 47048
rect 22704 46996 22710 47048
rect 13403 46971 13461 46977
rect 13403 46937 13415 46971
rect 13449 46968 13461 46971
rect 14274 46968 14280 46980
rect 13449 46940 14280 46968
rect 13449 46937 13461 46940
rect 13403 46931 13461 46937
rect 14274 46928 14280 46940
rect 14332 46928 14338 46980
rect 14458 46928 14464 46980
rect 14516 46928 14522 46980
rect 16117 46971 16175 46977
rect 16117 46937 16129 46971
rect 16163 46968 16175 46971
rect 20438 46968 20444 46980
rect 16163 46940 20444 46968
rect 16163 46937 16175 46940
rect 16117 46931 16175 46937
rect 20438 46928 20444 46940
rect 20496 46928 20502 46980
rect 20806 46928 20812 46980
rect 20864 46968 20870 46980
rect 23293 46971 23351 46977
rect 23293 46968 23305 46971
rect 20864 46940 23305 46968
rect 20864 46928 20870 46940
rect 23293 46937 23305 46940
rect 23339 46937 23351 46971
rect 23293 46931 23351 46937
rect 25314 46860 25320 46912
rect 25372 46900 25378 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 25372 46872 25421 46900
rect 25372 46860 25378 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 11422 46588 11428 46640
rect 11480 46628 11486 46640
rect 12345 46631 12403 46637
rect 12345 46628 12357 46631
rect 11480 46600 12357 46628
rect 11480 46588 11486 46600
rect 12345 46597 12357 46600
rect 12391 46597 12403 46631
rect 12345 46591 12403 46597
rect 14642 46588 14648 46640
rect 14700 46588 14706 46640
rect 25314 46520 25320 46572
rect 25372 46520 25378 46572
rect 12161 46495 12219 46501
rect 12161 46461 12173 46495
rect 12207 46492 12219 46495
rect 13538 46492 13544 46504
rect 12207 46464 13544 46492
rect 12207 46461 12219 46464
rect 12161 46455 12219 46461
rect 13538 46452 13544 46464
rect 13596 46452 13602 46504
rect 14001 46495 14059 46501
rect 14001 46461 14013 46495
rect 14047 46461 14059 46495
rect 14001 46455 14059 46461
rect 14461 46495 14519 46501
rect 14461 46461 14473 46495
rect 14507 46492 14519 46495
rect 15654 46492 15660 46504
rect 14507 46464 15660 46492
rect 14507 46461 14519 46464
rect 14461 46455 14519 46461
rect 14016 46424 14044 46455
rect 15654 46452 15660 46464
rect 15712 46452 15718 46504
rect 16301 46495 16359 46501
rect 16301 46461 16313 46495
rect 16347 46492 16359 46495
rect 21726 46492 21732 46504
rect 16347 46464 21732 46492
rect 16347 46461 16359 46464
rect 16301 46455 16359 46461
rect 21726 46452 21732 46464
rect 21784 46452 21790 46504
rect 19702 46424 19708 46436
rect 14016 46396 19708 46424
rect 19702 46384 19708 46396
rect 19760 46384 19766 46436
rect 22646 46316 22652 46368
rect 22704 46356 22710 46368
rect 25133 46359 25191 46365
rect 25133 46356 25145 46359
rect 22704 46328 25145 46356
rect 22704 46316 22710 46328
rect 25133 46325 25145 46328
rect 25179 46325 25191 46359
rect 25133 46319 25191 46325
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 9766 46112 9772 46164
rect 9824 46112 9830 46164
rect 10134 46016 10140 46028
rect 9140 45988 10140 46016
rect 9140 45957 9168 45988
rect 10134 45976 10140 45988
rect 10192 45976 10198 46028
rect 10778 45976 10784 46028
rect 10836 45976 10842 46028
rect 12066 45976 12072 46028
rect 12124 45976 12130 46028
rect 14274 45976 14280 46028
rect 14332 46016 14338 46028
rect 15749 46019 15807 46025
rect 15749 46016 15761 46019
rect 14332 45988 15761 46016
rect 14332 45976 14338 45988
rect 15749 45985 15761 45988
rect 15795 45985 15807 46019
rect 15749 45979 15807 45985
rect 9125 45951 9183 45957
rect 9125 45917 9137 45951
rect 9171 45917 9183 45951
rect 9125 45911 9183 45917
rect 9306 45908 9312 45960
rect 9364 45948 9370 45960
rect 10597 45951 10655 45957
rect 10597 45948 10609 45951
rect 9364 45920 10609 45948
rect 9364 45908 9370 45920
rect 10597 45917 10609 45920
rect 10643 45917 10655 45951
rect 10597 45911 10655 45917
rect 15565 45951 15623 45957
rect 15565 45917 15577 45951
rect 15611 45917 15623 45951
rect 15565 45911 15623 45917
rect 24857 45951 24915 45957
rect 24857 45917 24869 45951
rect 24903 45948 24915 45951
rect 25314 45948 25320 45960
rect 24903 45920 25320 45948
rect 24903 45917 24915 45920
rect 24857 45911 24915 45917
rect 15580 45812 15608 45911
rect 25314 45908 25320 45920
rect 25372 45908 25378 45960
rect 17126 45880 17132 45892
rect 16546 45852 17132 45880
rect 16546 45812 16574 45852
rect 17126 45840 17132 45852
rect 17184 45840 17190 45892
rect 17405 45883 17463 45889
rect 17405 45849 17417 45883
rect 17451 45880 17463 45883
rect 20162 45880 20168 45892
rect 17451 45852 20168 45880
rect 17451 45849 17463 45852
rect 17405 45843 17463 45849
rect 20162 45840 20168 45852
rect 20220 45840 20226 45892
rect 15580 45784 16574 45812
rect 22462 45772 22468 45824
rect 22520 45812 22526 45824
rect 25133 45815 25191 45821
rect 25133 45812 25145 45815
rect 22520 45784 25145 45812
rect 22520 45772 22526 45784
rect 25133 45781 25145 45784
rect 25179 45781 25191 45815
rect 25133 45775 25191 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 10778 45568 10784 45620
rect 10836 45608 10842 45620
rect 12158 45608 12164 45620
rect 10836 45580 12164 45608
rect 10836 45568 10842 45580
rect 12158 45568 12164 45580
rect 12216 45568 12222 45620
rect 9490 45500 9496 45552
rect 9548 45500 9554 45552
rect 11146 45432 11152 45484
rect 11204 45472 11210 45484
rect 11701 45475 11759 45481
rect 11701 45472 11713 45475
rect 11204 45444 11713 45472
rect 11204 45432 11210 45444
rect 11701 45441 11713 45444
rect 11747 45472 11759 45475
rect 12529 45475 12587 45481
rect 12529 45472 12541 45475
rect 11747 45444 12541 45472
rect 11747 45441 11759 45444
rect 11701 45435 11759 45441
rect 12529 45441 12541 45444
rect 12575 45441 12587 45475
rect 12529 45435 12587 45441
rect 9030 45364 9036 45416
rect 9088 45404 9094 45416
rect 9309 45407 9367 45413
rect 9309 45404 9321 45407
rect 9088 45376 9321 45404
rect 9088 45364 9094 45376
rect 9309 45373 9321 45376
rect 9355 45373 9367 45407
rect 9309 45367 9367 45373
rect 10962 45364 10968 45416
rect 11020 45364 11026 45416
rect 11790 45228 11796 45280
rect 11848 45228 11854 45280
rect 25314 45228 25320 45280
rect 25372 45268 25378 45280
rect 25409 45271 25467 45277
rect 25409 45268 25421 45271
rect 25372 45240 25421 45268
rect 25372 45228 25378 45240
rect 25409 45237 25421 45240
rect 25455 45237 25467 45271
rect 25409 45231 25467 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 10134 45024 10140 45076
rect 10192 45064 10198 45076
rect 10873 45067 10931 45073
rect 10873 45064 10885 45067
rect 10192 45036 10885 45064
rect 10192 45024 10198 45036
rect 10873 45033 10885 45036
rect 10919 45033 10931 45067
rect 10873 45027 10931 45033
rect 8570 44888 8576 44940
rect 8628 44928 8634 44940
rect 9125 44931 9183 44937
rect 9125 44928 9137 44931
rect 8628 44900 9137 44928
rect 8628 44888 8634 44900
rect 9125 44897 9137 44900
rect 9171 44928 9183 44931
rect 11514 44928 11520 44940
rect 9171 44900 11520 44928
rect 9171 44897 9183 44900
rect 9125 44891 9183 44897
rect 11514 44888 11520 44900
rect 11572 44888 11578 44940
rect 10502 44820 10508 44872
rect 10560 44820 10566 44872
rect 10870 44820 10876 44872
rect 10928 44860 10934 44872
rect 11333 44863 11391 44869
rect 11333 44860 11345 44863
rect 10928 44832 11345 44860
rect 10928 44820 10934 44832
rect 11333 44829 11345 44832
rect 11379 44829 11391 44863
rect 11333 44823 11391 44829
rect 25314 44820 25320 44872
rect 25372 44820 25378 44872
rect 9401 44795 9459 44801
rect 9401 44761 9413 44795
rect 9447 44761 9459 44795
rect 11977 44795 12035 44801
rect 11977 44792 11989 44795
rect 9401 44755 9459 44761
rect 10704 44764 11989 44792
rect 9416 44724 9444 44755
rect 10704 44724 10732 44764
rect 11977 44761 11989 44764
rect 12023 44761 12035 44795
rect 11977 44755 12035 44761
rect 9416 44696 10732 44724
rect 22370 44684 22376 44736
rect 22428 44724 22434 44736
rect 25133 44727 25191 44733
rect 25133 44724 25145 44727
rect 22428 44696 25145 44724
rect 22428 44684 22434 44696
rect 25133 44693 25145 44696
rect 25179 44693 25191 44727
rect 25133 44687 25191 44693
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 10870 44480 10876 44532
rect 10928 44480 10934 44532
rect 10226 44344 10232 44396
rect 10284 44344 10290 44396
rect 24762 44344 24768 44396
rect 24820 44384 24826 44396
rect 25133 44387 25191 44393
rect 25133 44384 25145 44387
rect 24820 44356 25145 44384
rect 24820 44344 24826 44356
rect 25133 44353 25145 44356
rect 25179 44353 25191 44387
rect 25133 44347 25191 44353
rect 11241 44319 11299 44325
rect 11241 44285 11253 44319
rect 11287 44316 11299 44319
rect 11514 44316 11520 44328
rect 11287 44288 11520 44316
rect 11287 44285 11299 44288
rect 11241 44279 11299 44285
rect 11514 44276 11520 44288
rect 11572 44276 11578 44328
rect 14366 44208 14372 44260
rect 14424 44248 14430 44260
rect 25317 44251 25375 44257
rect 25317 44248 25329 44251
rect 14424 44220 25329 44248
rect 14424 44208 14430 44220
rect 25317 44217 25329 44220
rect 25363 44217 25375 44251
rect 25317 44211 25375 44217
rect 10502 44140 10508 44192
rect 10560 44180 10566 44192
rect 11609 44183 11667 44189
rect 11609 44180 11621 44183
rect 10560 44152 11621 44180
rect 10560 44140 10566 44152
rect 11609 44149 11621 44152
rect 11655 44180 11667 44183
rect 11974 44180 11980 44192
rect 11655 44152 11980 44180
rect 11655 44149 11667 44152
rect 11609 44143 11667 44149
rect 11974 44140 11980 44152
rect 12032 44140 12038 44192
rect 19058 44140 19064 44192
rect 19116 44180 19122 44192
rect 25038 44180 25044 44192
rect 19116 44152 25044 44180
rect 19116 44140 19122 44152
rect 25038 44140 25044 44152
rect 25096 44140 25102 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 10226 43936 10232 43988
rect 10284 43976 10290 43988
rect 10597 43979 10655 43985
rect 10597 43976 10609 43979
rect 10284 43948 10609 43976
rect 10284 43936 10290 43948
rect 10597 43945 10609 43948
rect 10643 43945 10655 43979
rect 10597 43939 10655 43945
rect 20806 43800 20812 43852
rect 20864 43800 20870 43852
rect 21266 43800 21272 43852
rect 21324 43840 21330 43852
rect 22557 43843 22615 43849
rect 22557 43840 22569 43843
rect 21324 43812 22569 43840
rect 21324 43800 21330 43812
rect 22557 43809 22569 43812
rect 22603 43809 22615 43843
rect 22557 43803 22615 43809
rect 9950 43732 9956 43784
rect 10008 43772 10014 43784
rect 10318 43772 10324 43784
rect 10008 43744 10324 43772
rect 10008 43732 10014 43744
rect 10318 43732 10324 43744
rect 10376 43732 10382 43784
rect 19426 43732 19432 43784
rect 19484 43772 19490 43784
rect 20533 43775 20591 43781
rect 20533 43772 20545 43775
rect 19484 43744 20545 43772
rect 19484 43732 19490 43744
rect 20533 43741 20545 43744
rect 20579 43741 20591 43775
rect 20533 43735 20591 43741
rect 11974 43664 11980 43716
rect 12032 43704 12038 43716
rect 21082 43704 21088 43716
rect 12032 43676 21088 43704
rect 12032 43664 12038 43676
rect 21082 43664 21088 43676
rect 21140 43704 21146 43716
rect 21266 43704 21272 43716
rect 21140 43676 21272 43704
rect 21140 43664 21146 43676
rect 21266 43664 21272 43676
rect 21324 43664 21330 43716
rect 20622 43596 20628 43648
rect 20680 43636 20686 43648
rect 22281 43639 22339 43645
rect 22281 43636 22293 43639
rect 20680 43608 22293 43636
rect 20680 43596 20686 43608
rect 22281 43605 22293 43608
rect 22327 43605 22339 43639
rect 22281 43599 22339 43605
rect 25498 43596 25504 43648
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 25133 43367 25191 43373
rect 25133 43333 25145 43367
rect 25179 43364 25191 43367
rect 25498 43364 25504 43376
rect 25179 43336 25504 43364
rect 25179 43333 25191 43336
rect 25133 43327 25191 43333
rect 25498 43324 25504 43336
rect 25556 43324 25562 43376
rect 23474 43052 23480 43104
rect 23532 43092 23538 43104
rect 25225 43095 25283 43101
rect 25225 43092 25237 43095
rect 23532 43064 25237 43092
rect 23532 43052 23538 43064
rect 25225 43061 25237 43064
rect 25271 43061 25283 43095
rect 25225 43055 25283 43061
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 9940 42891 9998 42897
rect 9940 42857 9952 42891
rect 9986 42888 9998 42891
rect 11882 42888 11888 42900
rect 9986 42860 11888 42888
rect 9986 42857 9998 42860
rect 9940 42851 9998 42857
rect 11882 42848 11888 42860
rect 11940 42848 11946 42900
rect 9677 42755 9735 42761
rect 9677 42721 9689 42755
rect 9723 42752 9735 42755
rect 11514 42752 11520 42764
rect 9723 42724 11520 42752
rect 9723 42721 9735 42724
rect 9677 42715 9735 42721
rect 11514 42712 11520 42724
rect 11572 42712 11578 42764
rect 11974 42712 11980 42764
rect 12032 42712 12038 42764
rect 15930 42712 15936 42764
rect 15988 42752 15994 42764
rect 17310 42752 17316 42764
rect 15988 42724 17316 42752
rect 15988 42712 15994 42724
rect 17310 42712 17316 42724
rect 17368 42712 17374 42764
rect 11992 42684 12020 42712
rect 11086 42656 12020 42684
rect 24765 42619 24823 42625
rect 24765 42585 24777 42619
rect 24811 42616 24823 42619
rect 25130 42616 25136 42628
rect 24811 42588 25136 42616
rect 24811 42585 24823 42588
rect 24765 42579 24823 42585
rect 25130 42576 25136 42588
rect 25188 42576 25194 42628
rect 9950 42508 9956 42560
rect 10008 42548 10014 42560
rect 11425 42551 11483 42557
rect 11425 42548 11437 42551
rect 10008 42520 11437 42548
rect 10008 42508 10014 42520
rect 11425 42517 11437 42520
rect 11471 42517 11483 42551
rect 11425 42511 11483 42517
rect 11514 42508 11520 42560
rect 11572 42548 11578 42560
rect 11701 42551 11759 42557
rect 11701 42548 11713 42551
rect 11572 42520 11713 42548
rect 11572 42508 11578 42520
rect 11701 42517 11713 42520
rect 11747 42517 11759 42551
rect 11701 42511 11759 42517
rect 25222 42508 25228 42560
rect 25280 42508 25286 42560
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 25314 41964 25320 42016
rect 25372 42004 25378 42016
rect 25409 42007 25467 42013
rect 25409 42004 25421 42007
rect 25372 41976 25421 42004
rect 25372 41964 25378 41976
rect 25409 41973 25421 41976
rect 25455 41973 25467 42007
rect 25409 41967 25467 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 24765 41531 24823 41537
rect 24765 41497 24777 41531
rect 24811 41528 24823 41531
rect 25130 41528 25136 41540
rect 24811 41500 25136 41528
rect 24811 41497 24823 41500
rect 24765 41491 24823 41497
rect 25130 41488 25136 41500
rect 25188 41488 25194 41540
rect 16666 41420 16672 41472
rect 16724 41460 16730 41472
rect 23934 41460 23940 41472
rect 16724 41432 23940 41460
rect 16724 41420 16730 41432
rect 23934 41420 23940 41432
rect 23992 41420 23998 41472
rect 24854 41420 24860 41472
rect 24912 41460 24918 41472
rect 25225 41463 25283 41469
rect 25225 41460 25237 41463
rect 24912 41432 25237 41460
rect 24912 41420 24918 41432
rect 25225 41429 25237 41432
rect 25271 41429 25283 41463
rect 25225 41423 25283 41429
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 17218 41080 17224 41132
rect 17276 41120 17282 41132
rect 19429 41123 19487 41129
rect 19429 41120 19441 41123
rect 17276 41092 19441 41120
rect 17276 41080 17282 41092
rect 19429 41089 19441 41092
rect 19475 41120 19487 41123
rect 20622 41120 20628 41132
rect 19475 41092 20628 41120
rect 19475 41089 19487 41092
rect 19429 41083 19487 41089
rect 20622 41080 20628 41092
rect 20680 41080 20686 41132
rect 24213 41123 24271 41129
rect 24213 41089 24225 41123
rect 24259 41120 24271 41123
rect 24673 41123 24731 41129
rect 24673 41120 24685 41123
rect 24259 41092 24685 41120
rect 24259 41089 24271 41092
rect 24213 41083 24271 41089
rect 24673 41089 24685 41092
rect 24719 41120 24731 41123
rect 24854 41120 24860 41132
rect 24719 41092 24860 41120
rect 24719 41089 24731 41092
rect 24673 41083 24731 41089
rect 24854 41080 24860 41092
rect 24912 41080 24918 41132
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 18322 40876 18328 40928
rect 18380 40916 18386 40928
rect 20073 40919 20131 40925
rect 20073 40916 20085 40919
rect 18380 40888 20085 40916
rect 18380 40876 18386 40888
rect 20073 40885 20085 40888
rect 20119 40885 20131 40919
rect 20073 40879 20131 40885
rect 23842 40876 23848 40928
rect 23900 40916 23906 40928
rect 24489 40919 24547 40925
rect 24489 40916 24501 40919
rect 23900 40888 24501 40916
rect 23900 40876 23906 40888
rect 24489 40885 24501 40888
rect 24535 40885 24547 40919
rect 24489 40879 24547 40885
rect 24946 40876 24952 40928
rect 25004 40916 25010 40928
rect 25133 40919 25191 40925
rect 25133 40916 25145 40919
rect 25004 40888 25145 40916
rect 25004 40876 25010 40888
rect 25133 40885 25145 40888
rect 25179 40885 25191 40919
rect 25133 40879 25191 40885
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 25317 40511 25375 40517
rect 25317 40508 25329 40511
rect 24688 40480 25329 40508
rect 24688 40384 24716 40480
rect 25317 40477 25329 40480
rect 25363 40477 25375 40511
rect 25317 40471 25375 40477
rect 24670 40332 24676 40384
rect 24728 40332 24734 40384
rect 24762 40332 24768 40384
rect 24820 40372 24826 40384
rect 24857 40375 24915 40381
rect 24857 40372 24869 40375
rect 24820 40344 24869 40372
rect 24820 40332 24826 40344
rect 24857 40341 24869 40344
rect 24903 40341 24915 40375
rect 24857 40335 24915 40341
rect 25133 40375 25191 40381
rect 25133 40341 25145 40375
rect 25179 40372 25191 40375
rect 26142 40372 26148 40384
rect 25179 40344 26148 40372
rect 25179 40341 25191 40344
rect 25133 40335 25191 40341
rect 26142 40332 26148 40344
rect 26200 40332 26206 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 24762 40060 24768 40112
rect 24820 40100 24826 40112
rect 25133 40103 25191 40109
rect 25133 40100 25145 40103
rect 24820 40072 25145 40100
rect 24820 40060 24826 40072
rect 25133 40069 25145 40072
rect 25179 40069 25191 40103
rect 25133 40063 25191 40069
rect 24581 40035 24639 40041
rect 24581 40001 24593 40035
rect 24627 40032 24639 40035
rect 24854 40032 24860 40044
rect 24627 40004 24860 40032
rect 24627 40001 24639 40004
rect 24581 39995 24639 40001
rect 24854 39992 24860 40004
rect 24912 39992 24918 40044
rect 17034 39856 17040 39908
rect 17092 39896 17098 39908
rect 25317 39899 25375 39905
rect 25317 39896 25329 39899
rect 17092 39868 25329 39896
rect 17092 39856 17098 39868
rect 25317 39865 25329 39868
rect 25363 39865 25375 39899
rect 25317 39859 25375 39865
rect 24394 39788 24400 39840
rect 24452 39788 24458 39840
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 11882 39584 11888 39636
rect 11940 39584 11946 39636
rect 24765 39627 24823 39633
rect 24765 39593 24777 39627
rect 24811 39624 24823 39627
rect 24854 39624 24860 39636
rect 24811 39596 24860 39624
rect 24811 39593 24823 39596
rect 24765 39587 24823 39593
rect 24854 39584 24860 39596
rect 24912 39584 24918 39636
rect 11238 39380 11244 39432
rect 11296 39380 11302 39432
rect 24213 39355 24271 39361
rect 24213 39321 24225 39355
rect 24259 39352 24271 39355
rect 24302 39352 24308 39364
rect 24259 39324 24308 39352
rect 24259 39321 24271 39324
rect 24213 39315 24271 39321
rect 24302 39312 24308 39324
rect 24360 39352 24366 39364
rect 25133 39355 25191 39361
rect 25133 39352 25145 39355
rect 24360 39324 25145 39352
rect 24360 39312 24366 39324
rect 25133 39321 25145 39324
rect 25179 39321 25191 39355
rect 25133 39315 25191 39321
rect 25317 39355 25375 39361
rect 25317 39321 25329 39355
rect 25363 39352 25375 39355
rect 25498 39352 25504 39364
rect 25363 39324 25504 39352
rect 25363 39321 25375 39324
rect 25317 39315 25375 39321
rect 25498 39312 25504 39324
rect 25556 39312 25562 39364
rect 24486 39244 24492 39296
rect 24544 39244 24550 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 7742 39040 7748 39092
rect 7800 39080 7806 39092
rect 8573 39083 8631 39089
rect 8573 39080 8585 39083
rect 7800 39052 8585 39080
rect 7800 39040 7806 39052
rect 8573 39049 8585 39052
rect 8619 39049 8631 39083
rect 8573 39043 8631 39049
rect 8757 38947 8815 38953
rect 8757 38913 8769 38947
rect 8803 38944 8815 38947
rect 8846 38944 8852 38956
rect 8803 38916 8852 38944
rect 8803 38913 8815 38916
rect 8757 38907 8815 38913
rect 8846 38904 8852 38916
rect 8904 38904 8910 38956
rect 24213 38947 24271 38953
rect 24213 38913 24225 38947
rect 24259 38944 24271 38947
rect 24486 38944 24492 38956
rect 24259 38916 24492 38944
rect 24259 38913 24271 38916
rect 24213 38907 24271 38913
rect 24486 38904 24492 38916
rect 24544 38904 24550 38956
rect 24673 38947 24731 38953
rect 24673 38913 24685 38947
rect 24719 38944 24731 38947
rect 25130 38944 25136 38956
rect 24719 38916 25136 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 25130 38904 25136 38916
rect 25188 38904 25194 38956
rect 21082 38700 21088 38752
rect 21140 38740 21146 38752
rect 24029 38743 24087 38749
rect 24029 38740 24041 38743
rect 21140 38712 24041 38740
rect 21140 38700 21146 38712
rect 24029 38709 24041 38712
rect 24075 38709 24087 38743
rect 24029 38703 24087 38709
rect 25314 38700 25320 38752
rect 25372 38700 25378 38752
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 20070 38428 20076 38480
rect 20128 38468 20134 38480
rect 23845 38471 23903 38477
rect 23845 38468 23857 38471
rect 20128 38440 23857 38468
rect 20128 38428 20134 38440
rect 23845 38437 23857 38440
rect 23891 38437 23903 38471
rect 23845 38431 23903 38437
rect 18233 38335 18291 38341
rect 18233 38301 18245 38335
rect 18279 38332 18291 38335
rect 18322 38332 18328 38344
rect 18279 38304 18328 38332
rect 18279 38301 18291 38304
rect 18233 38295 18291 38301
rect 18322 38292 18328 38304
rect 18380 38292 18386 38344
rect 24029 38335 24087 38341
rect 24029 38332 24041 38335
rect 23492 38304 24041 38332
rect 14550 38156 14556 38208
rect 14608 38196 14614 38208
rect 18877 38199 18935 38205
rect 18877 38196 18889 38199
rect 14608 38168 18889 38196
rect 14608 38156 14614 38168
rect 18877 38165 18889 38168
rect 18923 38165 18935 38199
rect 18877 38159 18935 38165
rect 22738 38156 22744 38208
rect 22796 38196 22802 38208
rect 23492 38205 23520 38304
rect 24029 38301 24041 38304
rect 24075 38301 24087 38335
rect 24029 38295 24087 38301
rect 24578 38292 24584 38344
rect 24636 38292 24642 38344
rect 23477 38199 23535 38205
rect 23477 38196 23489 38199
rect 22796 38168 23489 38196
rect 22796 38156 22802 38168
rect 23477 38165 23489 38168
rect 23523 38165 23535 38199
rect 23477 38159 23535 38165
rect 24946 38156 24952 38208
rect 25004 38196 25010 38208
rect 25225 38199 25283 38205
rect 25225 38196 25237 38199
rect 25004 38168 25237 38196
rect 25004 38156 25010 38168
rect 25225 38165 25237 38168
rect 25271 38165 25283 38199
rect 25225 38159 25283 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 11238 37952 11244 38004
rect 11296 37992 11302 38004
rect 12345 37995 12403 38001
rect 12345 37992 12357 37995
rect 11296 37964 12357 37992
rect 11296 37952 11302 37964
rect 12345 37961 12357 37964
rect 12391 37961 12403 37995
rect 12345 37955 12403 37961
rect 11146 37816 11152 37868
rect 11204 37856 11210 37868
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 11204 37828 11713 37856
rect 11204 37816 11210 37828
rect 11701 37825 11713 37828
rect 11747 37856 11759 37859
rect 11790 37856 11796 37868
rect 11747 37828 11796 37856
rect 11747 37825 11759 37828
rect 11701 37819 11759 37825
rect 11790 37816 11796 37828
rect 11848 37816 11854 37868
rect 17310 37816 17316 37868
rect 17368 37856 17374 37868
rect 23017 37859 23075 37865
rect 23017 37856 23029 37859
rect 17368 37828 23029 37856
rect 17368 37816 17374 37828
rect 23017 37825 23029 37828
rect 23063 37825 23075 37859
rect 23017 37819 23075 37825
rect 23658 37816 23664 37868
rect 23716 37856 23722 37868
rect 24029 37859 24087 37865
rect 24029 37856 24041 37859
rect 23716 37828 24041 37856
rect 23716 37816 23722 37828
rect 24029 37825 24041 37828
rect 24075 37825 24087 37859
rect 24029 37819 24087 37825
rect 22741 37791 22799 37797
rect 22741 37757 22753 37791
rect 22787 37757 22799 37791
rect 22741 37751 22799 37757
rect 22756 37720 22784 37751
rect 24949 37723 25007 37729
rect 24949 37720 24961 37723
rect 22756 37692 24961 37720
rect 24949 37689 24961 37692
rect 24995 37720 25007 37723
rect 25038 37720 25044 37732
rect 24995 37692 25044 37720
rect 24995 37689 25007 37692
rect 24949 37683 25007 37689
rect 25038 37680 25044 37692
rect 25096 37680 25102 37732
rect 23474 37612 23480 37664
rect 23532 37652 23538 37664
rect 24673 37655 24731 37661
rect 24673 37652 24685 37655
rect 23532 37624 24685 37652
rect 23532 37612 23538 37624
rect 24673 37621 24685 37624
rect 24719 37621 24731 37655
rect 24673 37615 24731 37621
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 22281 37247 22339 37253
rect 22281 37213 22293 37247
rect 22327 37213 22339 37247
rect 22281 37207 22339 37213
rect 23385 37247 23443 37253
rect 23385 37213 23397 37247
rect 23431 37244 23443 37247
rect 23474 37244 23480 37256
rect 23431 37216 23480 37244
rect 23431 37213 23443 37216
rect 23385 37207 23443 37213
rect 22296 37176 22324 37207
rect 23474 37204 23480 37216
rect 23532 37204 23538 37256
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37244 24639 37247
rect 25222 37244 25228 37256
rect 24627 37216 25228 37244
rect 24627 37213 24639 37216
rect 24581 37207 24639 37213
rect 25222 37204 25228 37216
rect 25280 37204 25286 37256
rect 24029 37179 24087 37185
rect 24029 37176 24041 37179
rect 22296 37148 24041 37176
rect 24029 37145 24041 37148
rect 24075 37145 24087 37179
rect 24029 37139 24087 37145
rect 22186 37068 22192 37120
rect 22244 37108 22250 37120
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22244 37080 22937 37108
rect 22244 37068 22250 37080
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 22925 37071 22983 37077
rect 25225 37111 25283 37117
rect 25225 37077 25237 37111
rect 25271 37108 25283 37111
rect 25406 37108 25412 37120
rect 25271 37080 25412 37108
rect 25271 37077 25283 37080
rect 25225 37071 25283 37077
rect 25406 37068 25412 37080
rect 25464 37068 25470 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 20438 36864 20444 36916
rect 20496 36904 20502 36916
rect 20533 36907 20591 36913
rect 20533 36904 20545 36907
rect 20496 36876 20545 36904
rect 20496 36864 20502 36876
rect 20533 36873 20545 36876
rect 20579 36873 20591 36907
rect 20533 36867 20591 36873
rect 24213 36907 24271 36913
rect 24213 36873 24225 36907
rect 24259 36904 24271 36907
rect 24578 36904 24584 36916
rect 24259 36876 24584 36904
rect 24259 36873 24271 36876
rect 24213 36867 24271 36873
rect 24578 36864 24584 36876
rect 24636 36864 24642 36916
rect 25314 36836 25320 36848
rect 23584 36808 25320 36836
rect 22278 36728 22284 36780
rect 22336 36728 22342 36780
rect 23584 36777 23612 36808
rect 25314 36796 25320 36808
rect 25372 36796 25378 36848
rect 23569 36771 23627 36777
rect 23569 36737 23581 36771
rect 23615 36737 23627 36771
rect 23569 36731 23627 36737
rect 24673 36771 24731 36777
rect 24673 36737 24685 36771
rect 24719 36768 24731 36771
rect 24762 36768 24768 36780
rect 24719 36740 24768 36768
rect 24719 36737 24731 36740
rect 24673 36731 24731 36737
rect 24762 36728 24768 36740
rect 24820 36728 24826 36780
rect 22925 36567 22983 36573
rect 22925 36533 22937 36567
rect 22971 36564 22983 36567
rect 23382 36564 23388 36576
rect 22971 36536 23388 36564
rect 22971 36533 22983 36536
rect 22925 36527 22983 36533
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 24578 36524 24584 36576
rect 24636 36564 24642 36576
rect 25317 36567 25375 36573
rect 25317 36564 25329 36567
rect 24636 36536 25329 36564
rect 24636 36524 24642 36536
rect 25317 36533 25329 36536
rect 25363 36533 25375 36567
rect 25317 36527 25375 36533
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 22278 36320 22284 36372
rect 22336 36360 22342 36372
rect 23937 36363 23995 36369
rect 23937 36360 23949 36363
rect 22336 36332 23949 36360
rect 22336 36320 22342 36332
rect 23937 36329 23949 36332
rect 23983 36329 23995 36363
rect 23937 36323 23995 36329
rect 25222 36320 25228 36372
rect 25280 36320 25286 36372
rect 19978 36116 19984 36168
rect 20036 36116 20042 36168
rect 20625 36159 20683 36165
rect 20625 36125 20637 36159
rect 20671 36156 20683 36159
rect 21085 36159 21143 36165
rect 21085 36156 21097 36159
rect 20671 36128 21097 36156
rect 20671 36125 20683 36128
rect 20625 36119 20683 36125
rect 21085 36125 21097 36128
rect 21131 36125 21143 36159
rect 21085 36119 21143 36125
rect 21450 36116 21456 36168
rect 21508 36156 21514 36168
rect 22189 36159 22247 36165
rect 22189 36156 22201 36159
rect 21508 36128 22201 36156
rect 21508 36116 21514 36128
rect 22189 36125 22201 36128
rect 22235 36125 22247 36159
rect 22189 36119 22247 36125
rect 23290 36116 23296 36168
rect 23348 36116 23354 36168
rect 24578 36116 24584 36168
rect 24636 36116 24642 36168
rect 21729 36091 21787 36097
rect 21729 36057 21741 36091
rect 21775 36088 21787 36091
rect 24210 36088 24216 36100
rect 21775 36060 24216 36088
rect 21775 36057 21787 36060
rect 21729 36051 21787 36057
rect 24210 36048 24216 36060
rect 24268 36048 24274 36100
rect 22833 36023 22891 36029
rect 22833 35989 22845 36023
rect 22879 36020 22891 36023
rect 23198 36020 23204 36032
rect 22879 35992 23204 36020
rect 22879 35989 22891 35992
rect 22833 35983 22891 35989
rect 23198 35980 23204 35992
rect 23256 35980 23262 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 8754 35776 8760 35828
rect 8812 35776 8818 35828
rect 11514 35816 11520 35828
rect 9416 35788 11520 35816
rect 8941 35683 8999 35689
rect 8941 35649 8953 35683
rect 8987 35680 8999 35683
rect 9122 35680 9128 35692
rect 8987 35652 9128 35680
rect 8987 35649 8999 35652
rect 8941 35643 8999 35649
rect 9122 35640 9128 35652
rect 9180 35640 9186 35692
rect 9416 35689 9444 35788
rect 11514 35776 11520 35788
rect 11572 35776 11578 35828
rect 20438 35776 20444 35828
rect 20496 35816 20502 35828
rect 21085 35819 21143 35825
rect 21085 35816 21097 35819
rect 20496 35788 21097 35816
rect 20496 35776 20502 35788
rect 21085 35785 21097 35788
rect 21131 35785 21143 35819
rect 21085 35779 21143 35785
rect 11698 35748 11704 35760
rect 10902 35720 11704 35748
rect 11698 35708 11704 35720
rect 11756 35708 11762 35760
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35649 9459 35683
rect 9401 35643 9459 35649
rect 19150 35640 19156 35692
rect 19208 35680 19214 35692
rect 19613 35683 19671 35689
rect 19613 35680 19625 35683
rect 19208 35652 19625 35680
rect 19208 35640 19214 35652
rect 19613 35649 19625 35652
rect 19659 35649 19671 35683
rect 21100 35680 21128 35779
rect 22462 35776 22468 35828
rect 22520 35776 22526 35828
rect 21177 35751 21235 35757
rect 21177 35717 21189 35751
rect 21223 35748 21235 35751
rect 22646 35748 22652 35760
rect 21223 35720 22652 35748
rect 21223 35717 21235 35720
rect 21177 35711 21235 35717
rect 22646 35708 22652 35720
rect 22704 35708 22710 35760
rect 21100 35652 21404 35680
rect 19613 35643 19671 35649
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 11146 35572 11152 35624
rect 11204 35572 11210 35624
rect 21174 35572 21180 35624
rect 21232 35612 21238 35624
rect 21269 35615 21327 35621
rect 21269 35612 21281 35615
rect 21232 35584 21281 35612
rect 21232 35572 21238 35584
rect 21269 35581 21281 35584
rect 21315 35581 21327 35615
rect 21376 35612 21404 35652
rect 21726 35640 21732 35692
rect 21784 35680 21790 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 21784 35652 22385 35680
rect 21784 35640 21790 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 22480 35652 23152 35680
rect 22480 35612 22508 35652
rect 21376 35584 22508 35612
rect 21269 35575 21327 35581
rect 22554 35572 22560 35624
rect 22612 35572 22618 35624
rect 23124 35612 23152 35652
rect 23198 35640 23204 35692
rect 23256 35640 23262 35692
rect 23382 35640 23388 35692
rect 23440 35680 23446 35692
rect 24305 35683 24363 35689
rect 24305 35680 24317 35683
rect 23440 35652 24317 35680
rect 23440 35640 23446 35652
rect 24305 35649 24317 35652
rect 24351 35649 24363 35683
rect 24305 35643 24363 35649
rect 25866 35612 25872 35624
rect 23124 35584 25872 35612
rect 25866 35572 25872 35584
rect 25924 35572 25930 35624
rect 20806 35504 20812 35556
rect 20864 35544 20870 35556
rect 23845 35547 23903 35553
rect 23845 35544 23857 35547
rect 20864 35516 23857 35544
rect 20864 35504 20870 35516
rect 23845 35513 23857 35516
rect 23891 35513 23903 35547
rect 23845 35507 23903 35513
rect 11606 35436 11612 35488
rect 11664 35436 11670 35488
rect 20254 35436 20260 35488
rect 20312 35436 20318 35488
rect 20714 35436 20720 35488
rect 20772 35436 20778 35488
rect 20990 35436 20996 35488
rect 21048 35476 21054 35488
rect 22005 35479 22063 35485
rect 22005 35476 22017 35479
rect 21048 35448 22017 35476
rect 21048 35436 21054 35448
rect 22005 35445 22017 35448
rect 22051 35445 22063 35479
rect 22005 35439 22063 35445
rect 23934 35436 23940 35488
rect 23992 35476 23998 35488
rect 24949 35479 25007 35485
rect 24949 35476 24961 35479
rect 23992 35448 24961 35476
rect 23992 35436 23998 35448
rect 24949 35445 24961 35448
rect 24995 35445 25007 35479
rect 24949 35439 25007 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 18693 35275 18751 35281
rect 18693 35241 18705 35275
rect 18739 35272 18751 35275
rect 22278 35272 22284 35284
rect 18739 35244 22284 35272
rect 18739 35241 18751 35244
rect 18693 35235 18751 35241
rect 22278 35232 22284 35244
rect 22336 35232 22342 35284
rect 21726 35164 21732 35216
rect 21784 35164 21790 35216
rect 22097 35207 22155 35213
rect 22097 35173 22109 35207
rect 22143 35204 22155 35207
rect 22646 35204 22652 35216
rect 22143 35176 22652 35204
rect 22143 35173 22155 35176
rect 22097 35167 22155 35173
rect 22646 35164 22652 35176
rect 22704 35164 22710 35216
rect 19337 35139 19395 35145
rect 19337 35105 19349 35139
rect 19383 35136 19395 35139
rect 19383 35108 19417 35136
rect 19383 35105 19395 35108
rect 19337 35099 19395 35105
rect 18877 35071 18935 35077
rect 18877 35037 18889 35071
rect 18923 35068 18935 35071
rect 19352 35068 19380 35099
rect 20162 35096 20168 35148
rect 20220 35136 20226 35148
rect 20220 35108 22232 35136
rect 20220 35096 20226 35108
rect 18923 35040 19472 35068
rect 18923 35037 18935 35040
rect 18877 35031 18935 35037
rect 19444 35000 19472 35040
rect 19518 35028 19524 35080
rect 19576 35068 19582 35080
rect 19613 35071 19671 35077
rect 19613 35068 19625 35071
rect 19576 35040 19625 35068
rect 19576 35028 19582 35040
rect 19613 35037 19625 35040
rect 19659 35037 19671 35071
rect 19613 35031 19671 35037
rect 20254 35028 20260 35080
rect 20312 35068 20318 35080
rect 20717 35071 20775 35077
rect 20717 35068 20729 35071
rect 20312 35040 20729 35068
rect 20312 35028 20318 35040
rect 20717 35037 20729 35040
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 21818 35000 21824 35012
rect 19444 34972 21824 35000
rect 21818 34960 21824 34972
rect 21876 34960 21882 35012
rect 22204 35000 22232 35108
rect 22370 35096 22376 35148
rect 22428 35136 22434 35148
rect 23201 35139 23259 35145
rect 23201 35136 23213 35139
rect 22428 35108 23213 35136
rect 22428 35096 22434 35108
rect 23201 35105 23213 35108
rect 23247 35105 23259 35139
rect 23201 35099 23259 35105
rect 23290 35096 23296 35148
rect 23348 35096 23354 35148
rect 22281 35071 22339 35077
rect 22281 35037 22293 35071
rect 22327 35068 22339 35071
rect 23382 35068 23388 35080
rect 22327 35040 23388 35068
rect 22327 35037 22339 35040
rect 22281 35031 22339 35037
rect 23382 35028 23388 35040
rect 23440 35028 23446 35080
rect 24581 35071 24639 35077
rect 24581 35037 24593 35071
rect 24627 35068 24639 35071
rect 25222 35068 25228 35080
rect 24627 35040 25228 35068
rect 24627 35037 24639 35040
rect 24581 35031 24639 35037
rect 25222 35028 25228 35040
rect 25280 35028 25286 35080
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 22204 34972 23121 35000
rect 23109 34969 23121 34972
rect 23155 35000 23167 35003
rect 23937 35003 23995 35009
rect 23937 35000 23949 35003
rect 23155 34972 23949 35000
rect 23155 34969 23167 34972
rect 23109 34963 23167 34969
rect 23937 34969 23949 34972
rect 23983 35000 23995 35003
rect 24302 35000 24308 35012
rect 23983 34972 24308 35000
rect 23983 34969 23995 34972
rect 23937 34963 23995 34969
rect 24302 34960 24308 34972
rect 24360 34960 24366 35012
rect 18233 34935 18291 34941
rect 18233 34901 18245 34935
rect 18279 34932 18291 34935
rect 18322 34932 18328 34944
rect 18279 34904 18328 34932
rect 18279 34901 18291 34904
rect 18233 34895 18291 34901
rect 18322 34892 18328 34904
rect 18380 34892 18386 34944
rect 19610 34892 19616 34944
rect 19668 34932 19674 34944
rect 20257 34935 20315 34941
rect 20257 34932 20269 34935
rect 19668 34904 20269 34932
rect 19668 34892 19674 34904
rect 20257 34901 20269 34904
rect 20303 34901 20315 34935
rect 20257 34895 20315 34901
rect 20346 34892 20352 34944
rect 20404 34932 20410 34944
rect 21361 34935 21419 34941
rect 21361 34932 21373 34935
rect 20404 34904 21373 34932
rect 20404 34892 20410 34904
rect 21361 34901 21373 34904
rect 21407 34901 21419 34935
rect 21361 34895 21419 34901
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22520 34904 22753 34932
rect 22520 34892 22526 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 23753 34935 23811 34941
rect 23753 34932 23765 34935
rect 23440 34904 23765 34932
rect 23440 34892 23446 34904
rect 23753 34901 23765 34904
rect 23799 34901 23811 34935
rect 23753 34895 23811 34901
rect 24026 34892 24032 34944
rect 24084 34932 24090 34944
rect 24121 34935 24179 34941
rect 24121 34932 24133 34935
rect 24084 34904 24133 34932
rect 24084 34892 24090 34904
rect 24121 34901 24133 34904
rect 24167 34901 24179 34935
rect 24121 34895 24179 34901
rect 24946 34892 24952 34944
rect 25004 34932 25010 34944
rect 25225 34935 25283 34941
rect 25225 34932 25237 34935
rect 25004 34904 25237 34932
rect 25004 34892 25010 34904
rect 25225 34901 25237 34904
rect 25271 34901 25283 34935
rect 25225 34895 25283 34901
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 19150 34688 19156 34740
rect 19208 34688 19214 34740
rect 19702 34688 19708 34740
rect 19760 34728 19766 34740
rect 21361 34731 21419 34737
rect 21361 34728 21373 34731
rect 19760 34700 21373 34728
rect 19760 34688 19766 34700
rect 21361 34697 21373 34700
rect 21407 34697 21419 34731
rect 21361 34691 21419 34697
rect 21174 34660 21180 34672
rect 18524 34632 21180 34660
rect 18524 34601 18552 34632
rect 21174 34620 21180 34632
rect 21232 34620 21238 34672
rect 18049 34595 18107 34601
rect 18049 34561 18061 34595
rect 18095 34561 18107 34595
rect 18049 34555 18107 34561
rect 18509 34595 18567 34601
rect 18509 34561 18521 34595
rect 18555 34561 18567 34595
rect 18509 34555 18567 34561
rect 18064 34524 18092 34555
rect 19610 34552 19616 34604
rect 19668 34552 19674 34604
rect 20257 34595 20315 34601
rect 20257 34561 20269 34595
rect 20303 34592 20315 34595
rect 20717 34595 20775 34601
rect 20717 34592 20729 34595
rect 20303 34564 20729 34592
rect 20303 34561 20315 34564
rect 20257 34555 20315 34561
rect 20717 34561 20729 34564
rect 20763 34561 20775 34595
rect 20717 34555 20775 34561
rect 21358 34552 21364 34604
rect 21416 34592 21422 34604
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21416 34564 22017 34592
rect 21416 34552 21422 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22830 34552 22836 34604
rect 22888 34592 22894 34604
rect 23109 34595 23167 34601
rect 23109 34592 23121 34595
rect 22888 34564 23121 34592
rect 22888 34552 22894 34564
rect 23109 34561 23121 34564
rect 23155 34561 23167 34595
rect 23109 34555 23167 34561
rect 24210 34552 24216 34604
rect 24268 34552 24274 34604
rect 18322 34524 18328 34536
rect 18064 34496 18328 34524
rect 18322 34484 18328 34496
rect 18380 34524 18386 34536
rect 18380 34496 21588 34524
rect 18380 34484 18386 34496
rect 17034 34416 17040 34468
rect 17092 34456 17098 34468
rect 21560 34456 21588 34496
rect 22646 34484 22652 34536
rect 22704 34484 22710 34536
rect 23750 34484 23756 34536
rect 23808 34484 23814 34536
rect 24854 34484 24860 34536
rect 24912 34524 24918 34536
rect 25314 34524 25320 34536
rect 24912 34496 25320 34524
rect 24912 34484 24918 34496
rect 25314 34484 25320 34496
rect 25372 34484 25378 34536
rect 22094 34456 22100 34468
rect 17092 34428 21496 34456
rect 21560 34428 22100 34456
rect 17092 34416 17098 34428
rect 17865 34391 17923 34397
rect 17865 34357 17877 34391
rect 17911 34388 17923 34391
rect 19886 34388 19892 34400
rect 17911 34360 19892 34388
rect 17911 34357 17923 34360
rect 17865 34351 17923 34357
rect 19886 34348 19892 34360
rect 19944 34348 19950 34400
rect 21468 34388 21496 34428
rect 22094 34416 22100 34428
rect 22152 34416 22158 34468
rect 22554 34416 22560 34468
rect 22612 34416 22618 34468
rect 22572 34388 22600 34416
rect 23382 34388 23388 34400
rect 21468 34360 23388 34388
rect 23382 34348 23388 34360
rect 23440 34348 23446 34400
rect 24854 34348 24860 34400
rect 24912 34348 24918 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 9674 34144 9680 34196
rect 9732 34184 9738 34196
rect 10413 34187 10471 34193
rect 10413 34184 10425 34187
rect 9732 34156 10425 34184
rect 9732 34144 9738 34156
rect 10413 34153 10425 34156
rect 10459 34153 10471 34187
rect 10413 34147 10471 34153
rect 19692 34187 19750 34193
rect 19692 34153 19704 34187
rect 19738 34184 19750 34187
rect 24854 34184 24860 34196
rect 19738 34156 24860 34184
rect 19738 34153 19750 34156
rect 19692 34147 19750 34153
rect 24854 34144 24860 34156
rect 24912 34144 24918 34196
rect 25222 34144 25228 34196
rect 25280 34144 25286 34196
rect 21174 34076 21180 34128
rect 21232 34076 21238 34128
rect 23382 34076 23388 34128
rect 23440 34076 23446 34128
rect 11606 34008 11612 34060
rect 11664 34048 11670 34060
rect 15105 34051 15163 34057
rect 15105 34048 15117 34051
rect 11664 34020 15117 34048
rect 11664 34008 11670 34020
rect 15105 34017 15117 34020
rect 15151 34017 15163 34051
rect 15105 34011 15163 34017
rect 19426 34008 19432 34060
rect 19484 34048 19490 34060
rect 21634 34048 21640 34060
rect 19484 34020 21640 34048
rect 19484 34008 19490 34020
rect 21634 34008 21640 34020
rect 21692 34008 21698 34060
rect 9766 33940 9772 33992
rect 9824 33940 9830 33992
rect 17034 33940 17040 33992
rect 17092 33940 17098 33992
rect 18141 33983 18199 33989
rect 18141 33949 18153 33983
rect 18187 33980 18199 33983
rect 18322 33980 18328 33992
rect 18187 33952 18328 33980
rect 18187 33949 18199 33952
rect 18141 33943 18199 33949
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 24026 33940 24032 33992
rect 24084 33940 24090 33992
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33980 24639 33983
rect 25682 33980 25688 33992
rect 24627 33952 25688 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 25682 33940 25688 33952
rect 25740 33940 25746 33992
rect 14369 33915 14427 33921
rect 14369 33881 14381 33915
rect 14415 33912 14427 33915
rect 15378 33912 15384 33924
rect 14415 33884 15384 33912
rect 14415 33881 14427 33884
rect 14369 33875 14427 33881
rect 15378 33872 15384 33884
rect 15436 33912 15442 33924
rect 15565 33915 15623 33921
rect 15565 33912 15577 33915
rect 15436 33884 15577 33912
rect 15436 33872 15442 33884
rect 15565 33881 15577 33884
rect 15611 33881 15623 33915
rect 15565 33875 15623 33881
rect 17681 33915 17739 33921
rect 17681 33881 17693 33915
rect 17727 33912 17739 33915
rect 21174 33912 21180 33924
rect 17727 33884 19932 33912
rect 20930 33884 21180 33912
rect 17727 33881 17739 33884
rect 17681 33875 17739 33881
rect 18506 33804 18512 33856
rect 18564 33844 18570 33856
rect 18785 33847 18843 33853
rect 18785 33844 18797 33847
rect 18564 33816 18797 33844
rect 18564 33804 18570 33816
rect 18785 33813 18797 33816
rect 18831 33813 18843 33847
rect 19904 33844 19932 33884
rect 21174 33872 21180 33884
rect 21232 33872 21238 33924
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 22186 33912 22192 33924
rect 21959 33884 22192 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 22186 33872 22192 33884
rect 22244 33872 22250 33924
rect 22296 33884 22402 33912
rect 21450 33844 21456 33856
rect 19904 33816 21456 33844
rect 18785 33807 18843 33813
rect 21450 33804 21456 33816
rect 21508 33804 21514 33856
rect 22002 33804 22008 33856
rect 22060 33844 22066 33856
rect 22296 33844 22324 33884
rect 22060 33816 22324 33844
rect 23845 33847 23903 33853
rect 22060 33804 22066 33816
rect 23845 33813 23857 33847
rect 23891 33844 23903 33847
rect 25590 33844 25596 33856
rect 23891 33816 25596 33844
rect 23891 33813 23903 33816
rect 23845 33807 23903 33813
rect 25590 33804 25596 33816
rect 25648 33804 25654 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 16206 33600 16212 33652
rect 16264 33600 16270 33652
rect 16482 33600 16488 33652
rect 16540 33600 16546 33652
rect 18141 33643 18199 33649
rect 18141 33609 18153 33643
rect 18187 33640 18199 33643
rect 18322 33640 18328 33652
rect 18187 33612 18328 33640
rect 18187 33609 18199 33612
rect 18141 33603 18199 33609
rect 18322 33600 18328 33612
rect 18380 33600 18386 33652
rect 19978 33600 19984 33652
rect 20036 33640 20042 33652
rect 20438 33640 20444 33652
rect 20036 33612 20444 33640
rect 20036 33600 20042 33612
rect 20438 33600 20444 33612
rect 20496 33640 20502 33652
rect 21269 33643 21327 33649
rect 21269 33640 21281 33643
rect 20496 33612 21281 33640
rect 20496 33600 20502 33612
rect 21269 33609 21281 33612
rect 21315 33609 21327 33643
rect 22002 33640 22008 33652
rect 21269 33603 21327 33609
rect 21560 33612 22008 33640
rect 17497 33507 17555 33513
rect 17497 33473 17509 33507
rect 17543 33504 17555 33507
rect 18414 33504 18420 33516
rect 17543 33476 18420 33504
rect 17543 33473 17555 33476
rect 17497 33467 17555 33473
rect 18414 33464 18420 33476
rect 18472 33464 18478 33516
rect 18601 33507 18659 33513
rect 18601 33473 18613 33507
rect 18647 33504 18659 33507
rect 19061 33507 19119 33513
rect 19061 33504 19073 33507
rect 18647 33476 19073 33504
rect 18647 33473 18659 33476
rect 18601 33467 18659 33473
rect 19061 33473 19073 33476
rect 19107 33504 19119 33507
rect 19334 33504 19340 33516
rect 19107 33476 19340 33504
rect 19107 33473 19119 33476
rect 19061 33467 19119 33473
rect 19334 33464 19340 33476
rect 19392 33464 19398 33516
rect 20898 33464 20904 33516
rect 20956 33504 20962 33516
rect 21174 33504 21180 33516
rect 20956 33476 21180 33504
rect 20956 33464 20962 33476
rect 21174 33464 21180 33476
rect 21232 33504 21238 33516
rect 21560 33504 21588 33612
rect 22002 33600 22008 33612
rect 22060 33640 22066 33652
rect 22060 33612 22416 33640
rect 22060 33600 22066 33612
rect 21634 33532 21640 33584
rect 21692 33572 21698 33584
rect 22278 33572 22284 33584
rect 21692 33544 22284 33572
rect 21692 33532 21698 33544
rect 21232 33476 21588 33504
rect 21928 33504 21956 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 22388 33572 22416 33612
rect 23842 33600 23848 33652
rect 23900 33640 23906 33652
rect 24673 33643 24731 33649
rect 24673 33640 24685 33643
rect 23900 33612 24685 33640
rect 23900 33600 23906 33612
rect 24673 33609 24685 33612
rect 24719 33609 24731 33643
rect 24673 33603 24731 33609
rect 25222 33600 25228 33652
rect 25280 33640 25286 33652
rect 25317 33643 25375 33649
rect 25317 33640 25329 33643
rect 25280 33612 25329 33640
rect 25280 33600 25286 33612
rect 25317 33609 25329 33612
rect 25363 33640 25375 33643
rect 25866 33640 25872 33652
rect 25363 33612 25872 33640
rect 25363 33609 25375 33612
rect 25317 33603 25375 33609
rect 25866 33600 25872 33612
rect 25924 33600 25930 33652
rect 22388 33544 22770 33572
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21928 33476 22017 33504
rect 21232 33464 21238 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 24578 33464 24584 33516
rect 24636 33504 24642 33516
rect 25409 33507 25467 33513
rect 25409 33504 25421 33507
rect 24636 33476 25421 33504
rect 24636 33464 24642 33476
rect 25409 33473 25421 33476
rect 25455 33473 25467 33507
rect 25409 33467 25467 33473
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19521 33439 19579 33445
rect 19521 33436 19533 33439
rect 19484 33408 19533 33436
rect 19484 33396 19490 33408
rect 19521 33405 19533 33408
rect 19567 33405 19579 33439
rect 19521 33399 19579 33405
rect 19797 33439 19855 33445
rect 19797 33405 19809 33439
rect 19843 33436 19855 33439
rect 20806 33436 20812 33448
rect 19843 33408 20812 33436
rect 19843 33405 19855 33408
rect 19797 33399 19855 33405
rect 20806 33396 20812 33408
rect 20864 33396 20870 33448
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 23934 33436 23940 33448
rect 22327 33408 23940 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 24762 33396 24768 33448
rect 24820 33396 24826 33448
rect 18877 33303 18935 33309
rect 18877 33269 18889 33303
rect 18923 33300 18935 33303
rect 19242 33300 19248 33312
rect 18923 33272 19248 33300
rect 18923 33269 18935 33272
rect 18877 33263 18935 33269
rect 19242 33260 19248 33272
rect 19300 33260 19306 33312
rect 21637 33303 21695 33309
rect 21637 33269 21649 33303
rect 21683 33300 21695 33303
rect 22002 33300 22008 33312
rect 21683 33272 22008 33300
rect 21683 33269 21695 33272
rect 21637 33263 21695 33269
rect 22002 33260 22008 33272
rect 22060 33260 22066 33312
rect 23474 33260 23480 33312
rect 23532 33300 23538 33312
rect 23658 33300 23664 33312
rect 23532 33272 23664 33300
rect 23532 33260 23538 33272
rect 23658 33260 23664 33272
rect 23716 33300 23722 33312
rect 23753 33303 23811 33309
rect 23753 33300 23765 33303
rect 23716 33272 23765 33300
rect 23716 33260 23722 33272
rect 23753 33269 23765 33272
rect 23799 33269 23811 33303
rect 23753 33263 23811 33269
rect 24210 33260 24216 33312
rect 24268 33260 24274 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 9306 33056 9312 33108
rect 9364 33056 9370 33108
rect 18414 33056 18420 33108
rect 18472 33056 18478 33108
rect 18690 33056 18696 33108
rect 18748 33056 18754 33108
rect 18966 33056 18972 33108
rect 19024 33056 19030 33108
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 22094 33096 22100 33108
rect 19392 33068 22100 33096
rect 19392 33056 19398 33068
rect 22094 33056 22100 33068
rect 22152 33056 22158 33108
rect 22544 33099 22602 33105
rect 22544 33065 22556 33099
rect 22590 33096 22602 33099
rect 23198 33096 23204 33108
rect 22590 33068 23204 33096
rect 22590 33065 22602 33068
rect 22544 33059 22602 33065
rect 23198 33056 23204 33068
rect 23256 33056 23262 33108
rect 23290 33056 23296 33108
rect 23348 33096 23354 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 23348 33068 24041 33096
rect 23348 33056 23354 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 16025 32963 16083 32969
rect 16025 32929 16037 32963
rect 16071 32960 16083 32963
rect 17218 32960 17224 32972
rect 16071 32932 17224 32960
rect 16071 32929 16083 32932
rect 16025 32923 16083 32929
rect 17218 32920 17224 32932
rect 17276 32920 17282 32972
rect 18984 32960 19012 33056
rect 20898 32988 20904 33040
rect 20956 33028 20962 33040
rect 21177 33031 21235 33037
rect 21177 33028 21189 33031
rect 20956 33000 21189 33028
rect 20956 32988 20962 33000
rect 21177 32997 21189 33000
rect 21223 33028 21235 33031
rect 21358 33028 21364 33040
rect 21223 33000 21364 33028
rect 21223 32997 21235 33000
rect 21177 32991 21235 32997
rect 21358 32988 21364 33000
rect 21416 32988 21422 33040
rect 24320 33000 25176 33028
rect 17696 32932 19012 32960
rect 19705 32963 19763 32969
rect 7742 32852 7748 32904
rect 7800 32892 7806 32904
rect 9493 32895 9551 32901
rect 9493 32892 9505 32895
rect 7800 32864 9505 32892
rect 7800 32852 7806 32864
rect 9493 32861 9505 32864
rect 9539 32861 9551 32895
rect 9493 32855 9551 32861
rect 15749 32895 15807 32901
rect 15749 32861 15761 32895
rect 15795 32892 15807 32895
rect 16482 32892 16488 32904
rect 15795 32864 16488 32892
rect 15795 32861 15807 32864
rect 15749 32855 15807 32861
rect 16482 32852 16488 32864
rect 16540 32852 16546 32904
rect 16945 32895 17003 32901
rect 16945 32861 16957 32895
rect 16991 32892 17003 32895
rect 17586 32892 17592 32904
rect 16991 32864 17592 32892
rect 16991 32861 17003 32864
rect 16945 32855 17003 32861
rect 17586 32852 17592 32864
rect 17644 32892 17650 32904
rect 17696 32892 17724 32932
rect 19705 32929 19717 32963
rect 19751 32960 19763 32963
rect 20346 32960 20352 32972
rect 19751 32932 20352 32960
rect 19751 32929 19763 32932
rect 19705 32923 19763 32929
rect 20346 32920 20352 32932
rect 20404 32920 20410 32972
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 22922 32920 22928 32972
rect 22980 32960 22986 32972
rect 24320 32960 24348 33000
rect 22980 32932 24348 32960
rect 22980 32920 22986 32932
rect 24394 32920 24400 32972
rect 24452 32960 24458 32972
rect 25148 32969 25176 33000
rect 25041 32963 25099 32969
rect 25041 32960 25053 32963
rect 24452 32932 25053 32960
rect 24452 32920 24458 32932
rect 25041 32929 25053 32932
rect 25087 32929 25099 32963
rect 25041 32923 25099 32929
rect 25133 32963 25191 32969
rect 25133 32929 25145 32963
rect 25179 32929 25191 32963
rect 25133 32923 25191 32929
rect 17644 32864 17724 32892
rect 17773 32895 17831 32901
rect 17644 32852 17650 32864
rect 17773 32861 17785 32895
rect 17819 32892 17831 32895
rect 18782 32892 18788 32904
rect 17819 32864 18788 32892
rect 17819 32861 17831 32864
rect 17773 32855 17831 32861
rect 18782 32852 18788 32864
rect 18840 32852 18846 32904
rect 19426 32852 19432 32904
rect 19484 32852 19490 32904
rect 20806 32852 20812 32904
rect 20864 32892 20870 32904
rect 21821 32895 21879 32901
rect 20864 32864 21036 32892
rect 20864 32852 20870 32864
rect 15841 32827 15899 32833
rect 15841 32793 15853 32827
rect 15887 32824 15899 32827
rect 16206 32824 16212 32836
rect 15887 32796 16212 32824
rect 15887 32793 15899 32796
rect 15841 32787 15899 32793
rect 16206 32784 16212 32796
rect 16264 32824 16270 32836
rect 16850 32824 16856 32836
rect 16264 32796 16856 32824
rect 16264 32784 16270 32796
rect 16850 32784 16856 32796
rect 16908 32784 16914 32836
rect 17037 32827 17095 32833
rect 17037 32793 17049 32827
rect 17083 32824 17095 32827
rect 18598 32824 18604 32836
rect 17083 32796 18604 32824
rect 17083 32793 17095 32796
rect 17037 32787 17095 32793
rect 18598 32784 18604 32796
rect 18656 32784 18662 32836
rect 20088 32796 20194 32824
rect 14734 32716 14740 32768
rect 14792 32756 14798 32768
rect 15381 32759 15439 32765
rect 15381 32756 15393 32759
rect 14792 32728 15393 32756
rect 14792 32716 14798 32728
rect 15381 32725 15393 32728
rect 15427 32725 15439 32759
rect 15381 32719 15439 32725
rect 16574 32716 16580 32768
rect 16632 32716 16638 32768
rect 18414 32716 18420 32768
rect 18472 32756 18478 32768
rect 20088 32756 20116 32796
rect 20824 32756 20852 32852
rect 21008 32824 21036 32864
rect 21821 32861 21833 32895
rect 21867 32892 21879 32895
rect 22002 32892 22008 32904
rect 21867 32864 22008 32892
rect 21867 32861 21879 32864
rect 21821 32855 21879 32861
rect 22002 32852 22008 32864
rect 22060 32852 22066 32904
rect 24949 32895 25007 32901
rect 24949 32861 24961 32895
rect 24995 32892 25007 32895
rect 25222 32892 25228 32904
rect 24995 32864 25228 32892
rect 24995 32861 25007 32864
rect 24949 32855 25007 32861
rect 25222 32852 25228 32864
rect 25280 32852 25286 32904
rect 23014 32824 23020 32836
rect 21008 32796 23020 32824
rect 23014 32784 23020 32796
rect 23072 32784 23078 32836
rect 25038 32824 25044 32836
rect 23860 32796 25044 32824
rect 18472 32728 20852 32756
rect 18472 32716 18478 32728
rect 21634 32716 21640 32768
rect 21692 32716 21698 32768
rect 23198 32716 23204 32768
rect 23256 32756 23262 32768
rect 23860 32756 23888 32796
rect 25038 32784 25044 32796
rect 25096 32784 25102 32836
rect 23256 32728 23888 32756
rect 23256 32716 23262 32728
rect 23934 32716 23940 32768
rect 23992 32756 23998 32768
rect 24581 32759 24639 32765
rect 24581 32756 24593 32759
rect 23992 32728 24593 32756
rect 23992 32716 23998 32728
rect 24581 32725 24593 32728
rect 24627 32725 24639 32759
rect 24581 32719 24639 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 9030 32512 9036 32564
rect 9088 32512 9094 32564
rect 21269 32555 21327 32561
rect 16868 32524 19932 32552
rect 15378 32444 15384 32496
rect 15436 32484 15442 32496
rect 16868 32493 16896 32524
rect 16853 32487 16911 32493
rect 16853 32484 16865 32487
rect 15436 32456 16865 32484
rect 15436 32444 15442 32456
rect 16853 32453 16865 32456
rect 16899 32453 16911 32487
rect 16853 32447 16911 32453
rect 18414 32444 18420 32496
rect 18472 32444 18478 32496
rect 19904 32493 19932 32524
rect 21269 32521 21281 32555
rect 21315 32552 21327 32555
rect 25038 32552 25044 32564
rect 21315 32524 25044 32552
rect 21315 32521 21327 32524
rect 21269 32515 21327 32521
rect 25038 32512 25044 32524
rect 25096 32512 25102 32564
rect 19889 32487 19947 32493
rect 19889 32453 19901 32487
rect 19935 32484 19947 32487
rect 21450 32484 21456 32496
rect 19935 32456 21456 32484
rect 19935 32453 19947 32456
rect 19889 32447 19947 32453
rect 21450 32444 21456 32456
rect 21508 32484 21514 32496
rect 22005 32487 22063 32493
rect 22005 32484 22017 32487
rect 21508 32456 22017 32484
rect 21508 32444 21514 32456
rect 22005 32453 22017 32456
rect 22051 32453 22063 32487
rect 22005 32447 22063 32453
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22741 32487 22799 32493
rect 22741 32484 22753 32487
rect 22336 32456 22753 32484
rect 22336 32444 22342 32456
rect 22741 32453 22753 32456
rect 22787 32453 22799 32487
rect 22741 32447 22799 32453
rect 9214 32376 9220 32428
rect 9272 32376 9278 32428
rect 22756 32416 22784 32447
rect 23014 32444 23020 32496
rect 23072 32484 23078 32496
rect 23072 32456 24150 32484
rect 23072 32444 23078 32456
rect 23382 32416 23388 32428
rect 22756 32388 23388 32416
rect 23382 32376 23388 32388
rect 23440 32376 23446 32428
rect 14274 32308 14280 32360
rect 14332 32348 14338 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 14332 32320 16129 32348
rect 14332 32308 14338 32320
rect 16117 32317 16129 32320
rect 16163 32348 16175 32351
rect 17126 32348 17132 32360
rect 16163 32320 17132 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 17126 32308 17132 32320
rect 17184 32348 17190 32360
rect 17681 32351 17739 32357
rect 17681 32348 17693 32351
rect 17184 32320 17693 32348
rect 17184 32308 17190 32320
rect 17681 32317 17693 32320
rect 17727 32317 17739 32351
rect 17681 32311 17739 32317
rect 17957 32351 18015 32357
rect 17957 32317 17969 32351
rect 18003 32348 18015 32351
rect 18506 32348 18512 32360
rect 18003 32320 18512 32348
rect 18003 32317 18015 32320
rect 17957 32311 18015 32317
rect 18506 32308 18512 32320
rect 18564 32308 18570 32360
rect 19426 32308 19432 32360
rect 19484 32348 19490 32360
rect 20622 32348 20628 32360
rect 19484 32320 20628 32348
rect 19484 32308 19490 32320
rect 20622 32308 20628 32320
rect 20680 32308 20686 32360
rect 23661 32351 23719 32357
rect 23661 32317 23673 32351
rect 23707 32348 23719 32351
rect 25406 32348 25412 32360
rect 23707 32320 25412 32348
rect 23707 32317 23719 32320
rect 23661 32311 23719 32317
rect 25406 32308 25412 32320
rect 25464 32308 25470 32360
rect 15010 32172 15016 32224
rect 15068 32212 15074 32224
rect 16669 32215 16727 32221
rect 16669 32212 16681 32215
rect 15068 32184 16681 32212
rect 15068 32172 15074 32184
rect 16669 32181 16681 32184
rect 16715 32181 16727 32215
rect 16669 32175 16727 32181
rect 19429 32215 19487 32221
rect 19429 32181 19441 32215
rect 19475 32212 19487 32215
rect 19518 32212 19524 32224
rect 19475 32184 19524 32212
rect 19475 32181 19487 32184
rect 19429 32175 19487 32181
rect 19518 32172 19524 32184
rect 19576 32212 19582 32224
rect 22554 32212 22560 32224
rect 19576 32184 22560 32212
rect 19576 32172 19582 32184
rect 22554 32172 22560 32184
rect 22612 32172 22618 32224
rect 25130 32172 25136 32224
rect 25188 32172 25194 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 9766 31968 9772 32020
rect 9824 32008 9830 32020
rect 9861 32011 9919 32017
rect 9861 32008 9873 32011
rect 9824 31980 9873 32008
rect 9824 31968 9830 31980
rect 9861 31977 9873 31980
rect 9907 31977 9919 32011
rect 9861 31971 9919 31977
rect 13906 31968 13912 32020
rect 13964 32008 13970 32020
rect 16025 32011 16083 32017
rect 16025 32008 16037 32011
rect 13964 31980 16037 32008
rect 13964 31968 13970 31980
rect 16025 31977 16037 31980
rect 16071 31977 16083 32011
rect 16025 31971 16083 31977
rect 16666 31968 16672 32020
rect 16724 31968 16730 32020
rect 19426 32008 19432 32020
rect 17052 31980 19432 32008
rect 12066 31900 12072 31952
rect 12124 31940 12130 31952
rect 13541 31943 13599 31949
rect 13541 31940 13553 31943
rect 12124 31912 13553 31940
rect 12124 31900 12130 31912
rect 13541 31909 13553 31912
rect 13587 31909 13599 31943
rect 13541 31903 13599 31909
rect 16485 31943 16543 31949
rect 16485 31909 16497 31943
rect 16531 31940 16543 31943
rect 16942 31940 16948 31952
rect 16531 31912 16948 31940
rect 16531 31909 16543 31912
rect 16485 31903 16543 31909
rect 16942 31900 16948 31912
rect 17000 31900 17006 31952
rect 10502 31832 10508 31884
rect 10560 31872 10566 31884
rect 12345 31875 12403 31881
rect 12345 31872 12357 31875
rect 10560 31844 12357 31872
rect 10560 31832 10566 31844
rect 12345 31841 12357 31844
rect 12391 31841 12403 31875
rect 12345 31835 12403 31841
rect 12618 31832 12624 31884
rect 12676 31872 12682 31884
rect 14274 31872 14280 31884
rect 12676 31844 14280 31872
rect 12676 31832 12682 31844
rect 14274 31832 14280 31844
rect 14332 31832 14338 31884
rect 14550 31832 14556 31884
rect 14608 31832 14614 31884
rect 17052 31881 17080 31980
rect 19426 31968 19432 31980
rect 19484 31968 19490 32020
rect 20806 31968 20812 32020
rect 20864 32008 20870 32020
rect 21177 32011 21235 32017
rect 21177 32008 21189 32011
rect 20864 31980 21189 32008
rect 20864 31968 20870 31980
rect 21177 31977 21189 31980
rect 21223 31977 21235 32011
rect 21177 31971 21235 31977
rect 21450 31968 21456 32020
rect 21508 31968 21514 32020
rect 21634 31968 21640 32020
rect 21692 32008 21698 32020
rect 25406 32008 25412 32020
rect 21692 31980 25412 32008
rect 21692 31968 21698 31980
rect 25406 31968 25412 31980
rect 25464 31968 25470 32020
rect 18782 31900 18788 31952
rect 18840 31900 18846 31952
rect 23845 31943 23903 31949
rect 23845 31940 23857 31943
rect 19352 31912 19564 31940
rect 17037 31875 17095 31881
rect 17037 31841 17049 31875
rect 17083 31841 17095 31875
rect 17037 31835 17095 31841
rect 17313 31875 17371 31881
rect 17313 31841 17325 31875
rect 17359 31872 17371 31875
rect 19352 31872 19380 31912
rect 17359 31844 19380 31872
rect 19536 31872 19564 31912
rect 20732 31912 23857 31940
rect 20732 31872 20760 31912
rect 23845 31909 23857 31912
rect 23891 31909 23903 31943
rect 23845 31903 23903 31909
rect 24854 31900 24860 31952
rect 24912 31940 24918 31952
rect 25225 31943 25283 31949
rect 25225 31940 25237 31943
rect 24912 31912 25237 31940
rect 24912 31900 24918 31912
rect 25225 31909 25237 31912
rect 25271 31909 25283 31943
rect 25225 31903 25283 31909
rect 19536 31844 20760 31872
rect 21008 31844 21772 31872
rect 17359 31841 17371 31844
rect 17313 31835 17371 31841
rect 9217 31807 9275 31813
rect 9217 31773 9229 31807
rect 9263 31804 9275 31807
rect 9674 31804 9680 31816
rect 9263 31776 9680 31804
rect 9263 31773 9275 31776
rect 9217 31767 9275 31773
rect 9674 31764 9680 31776
rect 9732 31764 9738 31816
rect 11146 31764 11152 31816
rect 11204 31804 11210 31816
rect 11701 31807 11759 31813
rect 11701 31804 11713 31807
rect 11204 31776 11713 31804
rect 11204 31764 11210 31776
rect 11701 31773 11713 31776
rect 11747 31773 11759 31807
rect 11701 31767 11759 31773
rect 12897 31807 12955 31813
rect 12897 31773 12909 31807
rect 12943 31804 12955 31807
rect 13998 31804 14004 31816
rect 12943 31776 14004 31804
rect 12943 31773 12955 31776
rect 12897 31767 12955 31773
rect 13998 31764 14004 31776
rect 14056 31764 14062 31816
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 13538 31696 13544 31748
rect 13596 31736 13602 31748
rect 15010 31736 15016 31748
rect 13596 31708 15016 31736
rect 13596 31696 13602 31708
rect 15010 31696 15016 31708
rect 15068 31696 15074 31748
rect 18690 31736 18696 31748
rect 18538 31708 18696 31736
rect 18690 31696 18696 31708
rect 18748 31736 18754 31748
rect 18748 31708 19334 31736
rect 18748 31696 18754 31708
rect 19306 31668 19334 31708
rect 19702 31696 19708 31748
rect 19760 31696 19766 31748
rect 20088 31708 20194 31736
rect 20088 31668 20116 31708
rect 19306 31640 20116 31668
rect 20530 31628 20536 31680
rect 20588 31668 20594 31680
rect 21008 31668 21036 31844
rect 21634 31764 21640 31816
rect 21692 31764 21698 31816
rect 21744 31804 21772 31844
rect 21818 31832 21824 31884
rect 21876 31872 21882 31884
rect 21876 31844 22140 31872
rect 21876 31832 21882 31844
rect 21744 31776 22048 31804
rect 22020 31677 22048 31776
rect 20588 31640 21036 31668
rect 22005 31671 22063 31677
rect 20588 31628 20594 31640
rect 22005 31637 22017 31671
rect 22051 31637 22063 31671
rect 22112 31668 22140 31844
rect 22554 31832 22560 31884
rect 22612 31832 22618 31884
rect 25314 31872 25320 31884
rect 23124 31844 25320 31872
rect 22465 31807 22523 31813
rect 22465 31773 22477 31807
rect 22511 31804 22523 31807
rect 23124 31804 23152 31844
rect 25314 31832 25320 31844
rect 25372 31832 25378 31884
rect 22511 31776 23152 31804
rect 22511 31773 22523 31776
rect 22465 31767 22523 31773
rect 23198 31764 23204 31816
rect 23256 31764 23262 31816
rect 24581 31807 24639 31813
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 25222 31804 25228 31816
rect 24627 31776 25228 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 22373 31671 22431 31677
rect 22373 31668 22385 31671
rect 22112 31640 22385 31668
rect 22005 31631 22063 31637
rect 22373 31637 22385 31640
rect 22419 31668 22431 31671
rect 24762 31668 24768 31680
rect 22419 31640 24768 31668
rect 22419 31637 22431 31640
rect 22373 31631 22431 31637
rect 24762 31628 24768 31640
rect 24820 31628 24826 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 19702 31424 19708 31476
rect 19760 31464 19766 31476
rect 20162 31464 20168 31476
rect 19760 31436 20168 31464
rect 19760 31424 19766 31436
rect 20162 31424 20168 31436
rect 20220 31424 20226 31476
rect 20254 31424 20260 31476
rect 20312 31464 20318 31476
rect 20625 31467 20683 31473
rect 20625 31464 20637 31467
rect 20312 31436 20637 31464
rect 20312 31424 20318 31436
rect 20625 31433 20637 31436
rect 20671 31433 20683 31467
rect 20625 31427 20683 31433
rect 21450 31424 21456 31476
rect 21508 31464 21514 31476
rect 21545 31467 21603 31473
rect 21545 31464 21557 31467
rect 21508 31436 21557 31464
rect 21508 31424 21514 31436
rect 21545 31433 21557 31436
rect 21591 31433 21603 31467
rect 21545 31427 21603 31433
rect 22649 31467 22707 31473
rect 22649 31433 22661 31467
rect 22695 31464 22707 31467
rect 23198 31464 23204 31476
rect 22695 31436 23204 31464
rect 22695 31433 22707 31436
rect 22649 31427 22707 31433
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 24670 31424 24676 31476
rect 24728 31464 24734 31476
rect 25133 31467 25191 31473
rect 25133 31464 25145 31467
rect 24728 31436 25145 31464
rect 24728 31424 24734 31436
rect 25133 31433 25145 31436
rect 25179 31433 25191 31467
rect 25133 31427 25191 31433
rect 14001 31399 14059 31405
rect 14001 31396 14013 31399
rect 12268 31368 14013 31396
rect 10505 31331 10563 31337
rect 10505 31297 10517 31331
rect 10551 31328 10563 31331
rect 11238 31328 11244 31340
rect 10551 31300 11244 31328
rect 10551 31297 10563 31300
rect 10505 31291 10563 31297
rect 11238 31288 11244 31300
rect 11296 31288 11302 31340
rect 12268 31337 12296 31368
rect 14001 31365 14013 31368
rect 14047 31365 14059 31399
rect 17037 31399 17095 31405
rect 17037 31396 17049 31399
rect 14001 31359 14059 31365
rect 15672 31368 17049 31396
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31297 12311 31331
rect 12253 31291 12311 31297
rect 13357 31331 13415 31337
rect 13357 31297 13369 31331
rect 13403 31328 13415 31331
rect 13906 31328 13912 31340
rect 13403 31300 13912 31328
rect 13403 31297 13415 31300
rect 13357 31291 13415 31297
rect 13906 31288 13912 31300
rect 13964 31288 13970 31340
rect 14550 31288 14556 31340
rect 14608 31288 14614 31340
rect 15672 31337 15700 31368
rect 17037 31365 17049 31368
rect 17083 31396 17095 31399
rect 23934 31396 23940 31408
rect 17083 31368 23940 31396
rect 17083 31365 17095 31368
rect 17037 31359 17095 31365
rect 23934 31356 23940 31368
rect 23992 31356 23998 31408
rect 24118 31356 24124 31408
rect 24176 31356 24182 31408
rect 15657 31331 15715 31337
rect 15657 31297 15669 31331
rect 15703 31297 15715 31331
rect 15657 31291 15715 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31328 17371 31331
rect 17862 31328 17868 31340
rect 17359 31300 17868 31328
rect 17359 31297 17371 31300
rect 17313 31291 17371 31297
rect 17862 31288 17868 31300
rect 17920 31288 17926 31340
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31328 18015 31331
rect 18417 31331 18475 31337
rect 18417 31328 18429 31331
rect 18003 31300 18429 31328
rect 18003 31297 18015 31300
rect 17957 31291 18015 31297
rect 18417 31297 18429 31300
rect 18463 31297 18475 31331
rect 18417 31291 18475 31297
rect 20717 31331 20775 31337
rect 20717 31297 20729 31331
rect 20763 31328 20775 31331
rect 20763 31300 21404 31328
rect 20763 31297 20775 31300
rect 20717 31291 20775 31297
rect 19610 31220 19616 31272
rect 19668 31220 19674 31272
rect 19702 31220 19708 31272
rect 19760 31260 19766 31272
rect 20809 31263 20867 31269
rect 20809 31260 20821 31263
rect 19760 31232 20821 31260
rect 19760 31220 19766 31232
rect 20809 31229 20821 31232
rect 20855 31229 20867 31263
rect 21376 31260 21404 31300
rect 22002 31288 22008 31340
rect 22060 31288 22066 31340
rect 23382 31288 23388 31340
rect 23440 31288 23446 31340
rect 23661 31263 23719 31269
rect 21376 31232 22094 31260
rect 20809 31223 20867 31229
rect 10318 31152 10324 31204
rect 10376 31192 10382 31204
rect 12897 31195 12955 31201
rect 12897 31192 12909 31195
rect 10376 31164 12909 31192
rect 10376 31152 10382 31164
rect 12897 31161 12909 31164
rect 12943 31161 12955 31195
rect 12897 31155 12955 31161
rect 16301 31195 16359 31201
rect 16301 31161 16313 31195
rect 16347 31192 16359 31195
rect 21358 31192 21364 31204
rect 16347 31164 21364 31192
rect 16347 31161 16359 31164
rect 16301 31155 16359 31161
rect 21358 31152 21364 31164
rect 21416 31152 21422 31204
rect 9766 31084 9772 31136
rect 9824 31124 9830 31136
rect 11149 31127 11207 31133
rect 11149 31124 11161 31127
rect 9824 31096 11161 31124
rect 9824 31084 9830 31096
rect 11149 31093 11161 31096
rect 11195 31093 11207 31127
rect 11149 31087 11207 31093
rect 15197 31127 15255 31133
rect 15197 31093 15209 31127
rect 15243 31124 15255 31127
rect 16206 31124 16212 31136
rect 15243 31096 16212 31124
rect 15243 31093 15255 31096
rect 15197 31087 15255 31093
rect 16206 31084 16212 31096
rect 16264 31084 16270 31136
rect 16758 31084 16764 31136
rect 16816 31084 16822 31136
rect 17402 31084 17408 31136
rect 17460 31124 17466 31136
rect 19061 31127 19119 31133
rect 19061 31124 19073 31127
rect 17460 31096 19073 31124
rect 17460 31084 17466 31096
rect 19061 31093 19073 31096
rect 19107 31093 19119 31127
rect 19061 31087 19119 31093
rect 19518 31084 19524 31136
rect 19576 31124 19582 31136
rect 20257 31127 20315 31133
rect 20257 31124 20269 31127
rect 19576 31096 20269 31124
rect 19576 31084 19582 31096
rect 20257 31093 20269 31096
rect 20303 31093 20315 31127
rect 22066 31124 22094 31232
rect 23661 31229 23673 31263
rect 23707 31260 23719 31263
rect 24946 31260 24952 31272
rect 23707 31232 24952 31260
rect 23707 31229 23719 31232
rect 23661 31223 23719 31229
rect 24946 31220 24952 31232
rect 25004 31220 25010 31272
rect 26142 31124 26148 31136
rect 22066 31096 26148 31124
rect 20257 31087 20315 31093
rect 26142 31084 26148 31096
rect 26200 31084 26206 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 11238 30880 11244 30932
rect 11296 30880 11302 30932
rect 20254 30880 20260 30932
rect 20312 30920 20318 30932
rect 20349 30923 20407 30929
rect 20349 30920 20361 30923
rect 20312 30892 20361 30920
rect 20312 30880 20318 30892
rect 20349 30889 20361 30892
rect 20395 30889 20407 30923
rect 22002 30920 22008 30932
rect 20349 30883 20407 30889
rect 21008 30892 22008 30920
rect 15470 30812 15476 30864
rect 15528 30852 15534 30864
rect 15933 30855 15991 30861
rect 15933 30852 15945 30855
rect 15528 30824 15945 30852
rect 15528 30812 15534 30824
rect 15933 30821 15945 30824
rect 15979 30821 15991 30855
rect 15933 30815 15991 30821
rect 20073 30855 20131 30861
rect 20073 30821 20085 30855
rect 20119 30852 20131 30855
rect 21008 30852 21036 30892
rect 22002 30880 22008 30892
rect 22060 30880 22066 30932
rect 22830 30880 22836 30932
rect 22888 30880 22894 30932
rect 25222 30880 25228 30932
rect 25280 30880 25286 30932
rect 20119 30824 21036 30852
rect 20119 30821 20131 30824
rect 20073 30815 20131 30821
rect 23934 30812 23940 30864
rect 23992 30852 23998 30864
rect 25958 30852 25964 30864
rect 23992 30824 25964 30852
rect 23992 30812 23998 30824
rect 25958 30812 25964 30824
rect 26016 30812 26022 30864
rect 16482 30744 16488 30796
rect 16540 30744 16546 30796
rect 17126 30744 17132 30796
rect 17184 30744 17190 30796
rect 17402 30744 17408 30796
rect 17460 30744 17466 30796
rect 18877 30787 18935 30793
rect 18877 30753 18889 30787
rect 18923 30753 18935 30787
rect 18877 30747 18935 30753
rect 10134 30676 10140 30728
rect 10192 30716 10198 30728
rect 10597 30719 10655 30725
rect 10597 30716 10609 30719
rect 10192 30688 10609 30716
rect 10192 30676 10198 30688
rect 10597 30685 10609 30688
rect 10643 30685 10655 30719
rect 10597 30679 10655 30685
rect 11701 30719 11759 30725
rect 11701 30685 11713 30719
rect 11747 30685 11759 30719
rect 11701 30679 11759 30685
rect 11716 30648 11744 30679
rect 11790 30676 11796 30728
rect 11848 30716 11854 30728
rect 12805 30719 12863 30725
rect 12805 30716 12817 30719
rect 11848 30688 12817 30716
rect 11848 30676 11854 30688
rect 12805 30685 12817 30688
rect 12851 30685 12863 30719
rect 12805 30679 12863 30685
rect 15194 30676 15200 30728
rect 15252 30716 15258 30728
rect 16393 30719 16451 30725
rect 16393 30716 16405 30719
rect 15252 30688 16405 30716
rect 15252 30676 15258 30688
rect 16393 30685 16405 30688
rect 16439 30716 16451 30719
rect 16758 30716 16764 30728
rect 16439 30688 16764 30716
rect 16439 30685 16451 30688
rect 16393 30679 16451 30685
rect 16758 30676 16764 30688
rect 16816 30676 16822 30728
rect 18892 30716 18920 30747
rect 20622 30744 20628 30796
rect 20680 30784 20686 30796
rect 21085 30787 21143 30793
rect 21085 30784 21097 30787
rect 20680 30756 21097 30784
rect 20680 30744 20686 30756
rect 21085 30753 21097 30756
rect 21131 30753 21143 30787
rect 21085 30747 21143 30753
rect 21361 30787 21419 30793
rect 21361 30753 21373 30787
rect 21407 30784 21419 30787
rect 22830 30784 22836 30796
rect 21407 30756 22836 30784
rect 21407 30753 21419 30756
rect 21361 30747 21419 30753
rect 22830 30744 22836 30756
rect 22888 30744 22894 30796
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 18892 30688 19441 30716
rect 19429 30685 19441 30688
rect 19475 30716 19487 30719
rect 19702 30716 19708 30728
rect 19475 30688 19708 30716
rect 19475 30685 19487 30688
rect 19429 30679 19487 30685
rect 19702 30676 19708 30688
rect 19760 30676 19766 30728
rect 22646 30676 22652 30728
rect 22704 30716 22710 30728
rect 23293 30719 23351 30725
rect 23293 30716 23305 30719
rect 22704 30688 23305 30716
rect 22704 30676 22710 30688
rect 23293 30685 23305 30688
rect 23339 30685 23351 30719
rect 23293 30679 23351 30685
rect 24581 30719 24639 30725
rect 24581 30685 24593 30719
rect 24627 30685 24639 30719
rect 24581 30679 24639 30685
rect 12710 30648 12716 30660
rect 11716 30620 12716 30648
rect 12710 30608 12716 30620
rect 12768 30608 12774 30660
rect 14277 30651 14335 30657
rect 14277 30617 14289 30651
rect 14323 30617 14335 30651
rect 14277 30611 14335 30617
rect 11054 30540 11060 30592
rect 11112 30580 11118 30592
rect 12345 30583 12403 30589
rect 12345 30580 12357 30583
rect 11112 30552 12357 30580
rect 11112 30540 11118 30552
rect 12345 30549 12357 30552
rect 12391 30549 12403 30583
rect 12345 30543 12403 30549
rect 12894 30540 12900 30592
rect 12952 30580 12958 30592
rect 13449 30583 13507 30589
rect 13449 30580 13461 30583
rect 12952 30552 13461 30580
rect 12952 30540 12958 30552
rect 13449 30549 13461 30552
rect 13495 30549 13507 30583
rect 13449 30543 13507 30549
rect 13814 30540 13820 30592
rect 13872 30540 13878 30592
rect 14292 30580 14320 30611
rect 14366 30608 14372 30660
rect 14424 30648 14430 30660
rect 15013 30651 15071 30657
rect 15013 30648 15025 30651
rect 14424 30620 15025 30648
rect 14424 30608 14430 30620
rect 15013 30617 15025 30620
rect 15059 30617 15071 30651
rect 15013 30611 15071 30617
rect 15838 30608 15844 30660
rect 15896 30648 15902 30660
rect 16301 30651 16359 30657
rect 16301 30648 16313 30651
rect 15896 30620 16313 30648
rect 15896 30608 15902 30620
rect 16301 30617 16313 30620
rect 16347 30648 16359 30651
rect 16666 30648 16672 30660
rect 16347 30620 16672 30648
rect 16347 30617 16359 30620
rect 16301 30611 16359 30617
rect 16666 30608 16672 30620
rect 16724 30608 16730 30660
rect 18690 30648 18696 30660
rect 18630 30620 18696 30648
rect 18690 30608 18696 30620
rect 18748 30648 18754 30660
rect 21818 30648 21824 30660
rect 18748 30620 21824 30648
rect 18748 30608 18754 30620
rect 21818 30608 21824 30620
rect 21876 30608 21882 30660
rect 24596 30648 24624 30679
rect 23308 30620 24624 30648
rect 15378 30580 15384 30592
rect 14292 30552 15384 30580
rect 15378 30540 15384 30552
rect 15436 30580 15442 30592
rect 15565 30583 15623 30589
rect 15565 30580 15577 30583
rect 15436 30552 15577 30580
rect 15436 30540 15442 30552
rect 15565 30549 15577 30552
rect 15611 30580 15623 30583
rect 15746 30580 15752 30592
rect 15611 30552 15752 30580
rect 15611 30549 15623 30552
rect 15565 30543 15623 30549
rect 15746 30540 15752 30552
rect 15804 30540 15810 30592
rect 18414 30540 18420 30592
rect 18472 30580 18478 30592
rect 18708 30580 18736 30608
rect 18472 30552 18736 30580
rect 18472 30540 18478 30552
rect 20346 30540 20352 30592
rect 20404 30580 20410 30592
rect 20533 30583 20591 30589
rect 20533 30580 20545 30583
rect 20404 30552 20545 30580
rect 20404 30540 20410 30552
rect 20533 30549 20545 30552
rect 20579 30549 20591 30583
rect 20533 30543 20591 30549
rect 20806 30540 20812 30592
rect 20864 30580 20870 30592
rect 21174 30580 21180 30592
rect 20864 30552 21180 30580
rect 20864 30540 20870 30552
rect 21174 30540 21180 30552
rect 21232 30580 21238 30592
rect 23308 30580 23336 30620
rect 21232 30552 23336 30580
rect 23937 30583 23995 30589
rect 21232 30540 21238 30552
rect 23937 30549 23949 30583
rect 23983 30580 23995 30583
rect 24394 30580 24400 30592
rect 23983 30552 24400 30580
rect 23983 30549 23995 30552
rect 23937 30543 23995 30549
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 11698 30336 11704 30388
rect 11756 30376 11762 30388
rect 13538 30376 13544 30388
rect 11756 30348 13544 30376
rect 11756 30336 11762 30348
rect 9674 30268 9680 30320
rect 9732 30268 9738 30320
rect 11149 30311 11207 30317
rect 11149 30277 11161 30311
rect 11195 30308 11207 30311
rect 11790 30308 11796 30320
rect 11195 30280 11796 30308
rect 11195 30277 11207 30280
rect 11149 30271 11207 30277
rect 11790 30268 11796 30280
rect 11848 30268 11854 30320
rect 12894 30268 12900 30320
rect 12952 30268 12958 30320
rect 13359 30280 13387 30348
rect 13538 30336 13544 30348
rect 13596 30336 13602 30388
rect 14369 30379 14427 30385
rect 14369 30345 14381 30379
rect 14415 30376 14427 30379
rect 14550 30376 14556 30388
rect 14415 30348 14556 30376
rect 14415 30345 14427 30348
rect 14369 30339 14427 30345
rect 14550 30336 14556 30348
rect 14608 30376 14614 30388
rect 16482 30376 16488 30388
rect 14608 30348 16488 30376
rect 14608 30336 14614 30348
rect 16482 30336 16488 30348
rect 16540 30336 16546 30388
rect 17313 30379 17371 30385
rect 17313 30345 17325 30379
rect 17359 30345 17371 30379
rect 17313 30339 17371 30345
rect 16942 30268 16948 30320
rect 17000 30308 17006 30320
rect 17328 30308 17356 30339
rect 21818 30336 21824 30388
rect 21876 30376 21882 30388
rect 22278 30376 22284 30388
rect 21876 30348 22284 30376
rect 21876 30336 21882 30348
rect 22278 30336 22284 30348
rect 22336 30376 22342 30388
rect 22336 30348 24164 30376
rect 22336 30336 22342 30348
rect 17000 30280 17356 30308
rect 17000 30268 17006 30280
rect 17862 30268 17868 30320
rect 17920 30308 17926 30320
rect 18693 30311 18751 30317
rect 18693 30308 18705 30311
rect 17920 30280 18705 30308
rect 17920 30268 17926 30280
rect 18693 30277 18705 30280
rect 18739 30277 18751 30311
rect 18693 30271 18751 30277
rect 19058 30268 19064 30320
rect 19116 30308 19122 30320
rect 20162 30308 20168 30320
rect 19116 30280 20168 30308
rect 19116 30268 19122 30280
rect 20162 30268 20168 30280
rect 20220 30268 20226 30320
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 20990 30308 20996 30320
rect 20395 30280 20996 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 20990 30268 20996 30280
rect 21048 30268 21054 30320
rect 24136 30252 24164 30348
rect 9033 30243 9091 30249
rect 9033 30209 9045 30243
rect 9079 30240 9091 30243
rect 10226 30240 10232 30252
rect 9079 30212 10232 30240
rect 9079 30209 9091 30212
rect 9033 30203 9091 30209
rect 10226 30200 10232 30212
rect 10284 30200 10290 30252
rect 10502 30200 10508 30252
rect 10560 30200 10566 30252
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30240 14887 30243
rect 15746 30240 15752 30252
rect 14875 30212 15752 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 15746 30200 15752 30212
rect 15804 30200 15810 30252
rect 16298 30200 16304 30252
rect 16356 30240 16362 30252
rect 16393 30243 16451 30249
rect 16393 30240 16405 30243
rect 16356 30212 16405 30240
rect 16356 30200 16362 30212
rect 16393 30209 16405 30212
rect 16439 30209 16451 30243
rect 16393 30203 16451 30209
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 17221 30243 17279 30249
rect 16540 30212 17172 30240
rect 16540 30200 16546 30212
rect 12618 30132 12624 30184
rect 12676 30132 12682 30184
rect 14182 30132 14188 30184
rect 14240 30172 14246 30184
rect 15565 30175 15623 30181
rect 15565 30172 15577 30175
rect 14240 30144 15577 30172
rect 14240 30132 14246 30144
rect 15565 30141 15577 30144
rect 15611 30172 15623 30175
rect 17034 30172 17040 30184
rect 15611 30144 17040 30172
rect 15611 30141 15623 30144
rect 15565 30135 15623 30141
rect 17034 30132 17040 30144
rect 17092 30132 17098 30184
rect 17144 30172 17172 30212
rect 17221 30209 17233 30243
rect 17267 30240 17279 30243
rect 18049 30243 18107 30249
rect 17267 30212 17540 30240
rect 17267 30209 17279 30212
rect 17221 30203 17279 30209
rect 17405 30175 17463 30181
rect 17405 30172 17417 30175
rect 17144 30144 17417 30172
rect 17405 30141 17417 30144
rect 17451 30141 17463 30175
rect 17405 30135 17463 30141
rect 15746 30064 15752 30116
rect 15804 30104 15810 30116
rect 16301 30107 16359 30113
rect 16301 30104 16313 30107
rect 15804 30076 16313 30104
rect 15804 30064 15810 30076
rect 16301 30073 16313 30076
rect 16347 30104 16359 30107
rect 17218 30104 17224 30116
rect 16347 30076 17224 30104
rect 16347 30073 16359 30076
rect 16301 30067 16359 30073
rect 17218 30064 17224 30076
rect 17276 30064 17282 30116
rect 17512 30048 17540 30212
rect 18049 30209 18061 30243
rect 18095 30240 18107 30243
rect 18874 30240 18880 30252
rect 18095 30212 18880 30240
rect 18095 30209 18107 30212
rect 18049 30203 18107 30209
rect 18874 30200 18880 30212
rect 18932 30200 18938 30252
rect 18966 30200 18972 30252
rect 19024 30200 19030 30252
rect 19610 30200 19616 30252
rect 19668 30240 19674 30252
rect 20257 30243 20315 30249
rect 19668 30212 19932 30240
rect 19668 30200 19674 30212
rect 18322 30132 18328 30184
rect 18380 30172 18386 30184
rect 18984 30172 19012 30200
rect 18380 30144 19012 30172
rect 19153 30175 19211 30181
rect 18380 30132 18386 30144
rect 19153 30141 19165 30175
rect 19199 30172 19211 30175
rect 19794 30172 19800 30184
rect 19199 30144 19800 30172
rect 19199 30141 19211 30144
rect 19153 30135 19211 30141
rect 19794 30132 19800 30144
rect 19852 30132 19858 30184
rect 19904 30172 19932 30212
rect 20257 30209 20269 30243
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 21177 30243 21235 30249
rect 21177 30209 21189 30243
rect 21223 30209 21235 30243
rect 21177 30203 21235 30209
rect 22097 30243 22155 30249
rect 22097 30209 22109 30243
rect 22143 30209 22155 30243
rect 22097 30203 22155 30209
rect 20272 30172 20300 30203
rect 19904 30144 20300 30172
rect 20438 30132 20444 30184
rect 20496 30132 20502 30184
rect 18966 30064 18972 30116
rect 19024 30104 19030 30116
rect 21192 30104 21220 30203
rect 19024 30076 21220 30104
rect 21361 30107 21419 30113
rect 19024 30064 19030 30076
rect 21361 30073 21373 30107
rect 21407 30104 21419 30107
rect 21726 30104 21732 30116
rect 21407 30076 21732 30104
rect 21407 30073 21419 30076
rect 21361 30067 21419 30073
rect 21726 30064 21732 30076
rect 21784 30064 21790 30116
rect 15562 29996 15568 30048
rect 15620 30036 15626 30048
rect 16025 30039 16083 30045
rect 16025 30036 16037 30039
rect 15620 30008 16037 30036
rect 15620 29996 15626 30008
rect 16025 30005 16037 30008
rect 16071 30005 16083 30039
rect 16025 29999 16083 30005
rect 16758 29996 16764 30048
rect 16816 30036 16822 30048
rect 16853 30039 16911 30045
rect 16853 30036 16865 30039
rect 16816 30008 16865 30036
rect 16816 29996 16822 30008
rect 16853 30005 16865 30008
rect 16899 30005 16911 30039
rect 16853 29999 16911 30005
rect 17494 29996 17500 30048
rect 17552 30036 17558 30048
rect 19150 30036 19156 30048
rect 17552 30008 19156 30036
rect 17552 29996 17558 30008
rect 19150 29996 19156 30008
rect 19208 29996 19214 30048
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19889 30039 19947 30045
rect 19889 30036 19901 30039
rect 19392 30008 19901 30036
rect 19392 29996 19398 30008
rect 19889 30005 19901 30008
rect 19935 30005 19947 30039
rect 19889 29999 19947 30005
rect 20162 29996 20168 30048
rect 20220 30036 20226 30048
rect 22112 30036 22140 30203
rect 24118 30200 24124 30252
rect 24176 30200 24182 30252
rect 22738 30132 22744 30184
rect 22796 30132 22802 30184
rect 23017 30175 23075 30181
rect 23017 30141 23029 30175
rect 23063 30172 23075 30175
rect 23658 30172 23664 30184
rect 23063 30144 23664 30172
rect 23063 30141 23075 30144
rect 23017 30135 23075 30141
rect 23658 30132 23664 30144
rect 23716 30132 23722 30184
rect 24946 30132 24952 30184
rect 25004 30132 25010 30184
rect 22281 30107 22339 30113
rect 22281 30073 22293 30107
rect 22327 30104 22339 30107
rect 22554 30104 22560 30116
rect 22327 30076 22560 30104
rect 22327 30073 22339 30076
rect 22281 30067 22339 30073
rect 22554 30064 22560 30076
rect 22612 30064 22618 30116
rect 20220 30008 22140 30036
rect 20220 29996 20226 30008
rect 24486 29996 24492 30048
rect 24544 29996 24550 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 13814 29792 13820 29844
rect 13872 29832 13878 29844
rect 23382 29832 23388 29844
rect 13872 29804 23388 29832
rect 13872 29792 13878 29804
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 18506 29724 18512 29776
rect 18564 29764 18570 29776
rect 19334 29764 19340 29776
rect 18564 29736 19340 29764
rect 18564 29724 18570 29736
rect 19334 29724 19340 29736
rect 19392 29724 19398 29776
rect 20346 29724 20352 29776
rect 20404 29764 20410 29776
rect 20404 29736 21312 29764
rect 20404 29724 20410 29736
rect 11054 29696 11060 29708
rect 10152 29668 11060 29696
rect 10152 29637 10180 29668
rect 11054 29656 11060 29668
rect 11112 29656 11118 29708
rect 12526 29696 12532 29708
rect 11256 29668 12532 29696
rect 10137 29631 10195 29637
rect 10137 29597 10149 29631
rect 10183 29597 10195 29631
rect 10137 29591 10195 29597
rect 10870 29588 10876 29640
rect 10928 29628 10934 29640
rect 11256 29637 11284 29668
rect 12526 29656 12532 29668
rect 12584 29696 12590 29708
rect 14182 29696 14188 29708
rect 12584 29668 14188 29696
rect 12584 29656 12590 29668
rect 14182 29656 14188 29668
rect 14240 29656 14246 29708
rect 15286 29656 15292 29708
rect 15344 29696 15350 29708
rect 15565 29699 15623 29705
rect 15565 29696 15577 29699
rect 15344 29668 15577 29696
rect 15344 29656 15350 29668
rect 15565 29665 15577 29668
rect 15611 29696 15623 29699
rect 16114 29696 16120 29708
rect 15611 29668 16120 29696
rect 15611 29665 15623 29668
rect 15565 29659 15623 29665
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 16485 29699 16543 29705
rect 16485 29665 16497 29699
rect 16531 29696 16543 29699
rect 16850 29696 16856 29708
rect 16531 29668 16856 29696
rect 16531 29665 16543 29668
rect 16485 29659 16543 29665
rect 16850 29656 16856 29668
rect 16908 29656 16914 29708
rect 16942 29656 16948 29708
rect 17000 29696 17006 29708
rect 19150 29696 19156 29708
rect 17000 29668 19156 29696
rect 17000 29656 17006 29668
rect 19150 29656 19156 29668
rect 19208 29656 19214 29708
rect 20073 29699 20131 29705
rect 20073 29665 20085 29699
rect 20119 29696 20131 29699
rect 20898 29696 20904 29708
rect 20119 29668 20904 29696
rect 20119 29665 20131 29668
rect 20073 29659 20131 29665
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 11241 29631 11299 29637
rect 11241 29628 11253 29631
rect 10928 29600 11253 29628
rect 10928 29588 10934 29600
rect 11241 29597 11253 29600
rect 11287 29597 11299 29631
rect 11241 29591 11299 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 13814 29628 13820 29640
rect 13771 29600 13820 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 13814 29588 13820 29600
rect 13872 29588 13878 29640
rect 14553 29631 14611 29637
rect 14553 29597 14565 29631
rect 14599 29597 14611 29631
rect 14553 29591 14611 29597
rect 11514 29520 11520 29572
rect 11572 29520 11578 29572
rect 11790 29520 11796 29572
rect 11848 29560 11854 29572
rect 14568 29560 14596 29591
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 15381 29631 15439 29637
rect 15381 29628 15393 29631
rect 15068 29600 15393 29628
rect 15068 29588 15074 29600
rect 15381 29597 15393 29600
rect 15427 29628 15439 29631
rect 16298 29628 16304 29640
rect 15427 29600 16304 29628
rect 15427 29597 15439 29600
rect 15381 29591 15439 29597
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 17126 29588 17132 29640
rect 17184 29588 17190 29640
rect 19794 29588 19800 29640
rect 19852 29588 19858 29640
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29628 19947 29631
rect 20714 29628 20720 29640
rect 19935 29600 20720 29628
rect 19935 29597 19947 29600
rect 19889 29591 19947 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 21008 29637 21036 29736
rect 21082 29656 21088 29708
rect 21140 29656 21146 29708
rect 21177 29699 21235 29705
rect 21177 29665 21189 29699
rect 21223 29665 21235 29699
rect 21177 29659 21235 29665
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 16117 29563 16175 29569
rect 16117 29560 16129 29563
rect 11848 29532 12006 29560
rect 14568 29532 16129 29560
rect 11848 29520 11854 29532
rect 16117 29529 16129 29532
rect 16163 29560 16175 29563
rect 17310 29560 17316 29572
rect 16163 29532 17316 29560
rect 16163 29529 16175 29532
rect 16117 29523 16175 29529
rect 17310 29520 17316 29532
rect 17368 29520 17374 29572
rect 17402 29520 17408 29572
rect 17460 29520 17466 29572
rect 18414 29520 18420 29572
rect 18472 29520 18478 29572
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 21192 29560 21220 29659
rect 19392 29532 21220 29560
rect 19392 29520 19398 29532
rect 10781 29495 10839 29501
rect 10781 29461 10793 29495
rect 10827 29492 10839 29495
rect 11882 29492 11888 29504
rect 10827 29464 11888 29492
rect 10827 29461 10839 29464
rect 10781 29455 10839 29461
rect 11882 29452 11888 29464
rect 11940 29452 11946 29504
rect 12986 29452 12992 29504
rect 13044 29452 13050 29504
rect 13538 29452 13544 29504
rect 13596 29452 13602 29504
rect 14369 29495 14427 29501
rect 14369 29461 14381 29495
rect 14415 29492 14427 29495
rect 14550 29492 14556 29504
rect 14415 29464 14556 29492
rect 14415 29461 14427 29464
rect 14369 29455 14427 29461
rect 14550 29452 14556 29464
rect 14608 29452 14614 29504
rect 15013 29495 15071 29501
rect 15013 29461 15025 29495
rect 15059 29492 15071 29495
rect 15286 29492 15292 29504
rect 15059 29464 15292 29492
rect 15059 29461 15071 29464
rect 15013 29455 15071 29461
rect 15286 29452 15292 29464
rect 15344 29452 15350 29504
rect 15473 29495 15531 29501
rect 15473 29461 15485 29495
rect 15519 29492 15531 29495
rect 15746 29492 15752 29504
rect 15519 29464 15752 29492
rect 15519 29461 15531 29464
rect 15473 29455 15531 29461
rect 15746 29452 15752 29464
rect 15804 29452 15810 29504
rect 15930 29452 15936 29504
rect 15988 29492 15994 29504
rect 16298 29492 16304 29504
rect 15988 29464 16304 29492
rect 15988 29452 15994 29464
rect 16298 29452 16304 29464
rect 16356 29492 16362 29504
rect 18322 29492 18328 29504
rect 16356 29464 18328 29492
rect 16356 29452 16362 29464
rect 18322 29452 18328 29464
rect 18380 29452 18386 29504
rect 18874 29452 18880 29504
rect 18932 29452 18938 29504
rect 19429 29495 19487 29501
rect 19429 29461 19441 29495
rect 19475 29492 19487 29495
rect 19610 29492 19616 29504
rect 19475 29464 19616 29492
rect 19475 29461 19487 29464
rect 19429 29455 19487 29461
rect 19610 29452 19616 29464
rect 19668 29452 19674 29504
rect 20622 29452 20628 29504
rect 20680 29452 20686 29504
rect 21284 29492 21312 29736
rect 22830 29724 22836 29776
rect 22888 29764 22894 29776
rect 23937 29767 23995 29773
rect 23937 29764 23949 29767
rect 22888 29736 23949 29764
rect 22888 29724 22894 29736
rect 23937 29733 23949 29736
rect 23983 29733 23995 29767
rect 23937 29727 23995 29733
rect 24854 29696 24860 29708
rect 23308 29668 24860 29696
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 21910 29628 21916 29640
rect 21508 29600 21916 29628
rect 21508 29588 21514 29600
rect 21910 29588 21916 29600
rect 21968 29588 21974 29640
rect 23308 29637 23336 29668
rect 24854 29656 24860 29668
rect 24912 29656 24918 29708
rect 23293 29631 23351 29637
rect 23293 29597 23305 29631
rect 23339 29597 23351 29631
rect 23293 29591 23351 29597
rect 23750 29588 23756 29640
rect 23808 29628 23814 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 23808 29600 24593 29628
rect 23808 29588 23814 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 22094 29520 22100 29572
rect 22152 29560 22158 29572
rect 22649 29563 22707 29569
rect 22649 29560 22661 29563
rect 22152 29532 22661 29560
rect 22152 29520 22158 29532
rect 22649 29529 22661 29532
rect 22695 29560 22707 29563
rect 22738 29560 22744 29572
rect 22695 29532 22744 29560
rect 22695 29529 22707 29532
rect 22649 29523 22707 29529
rect 22738 29520 22744 29532
rect 22796 29520 22802 29572
rect 23566 29492 23572 29504
rect 21284 29464 23572 29492
rect 23566 29452 23572 29464
rect 23624 29452 23630 29504
rect 25222 29452 25228 29504
rect 25280 29452 25286 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 11514 29248 11520 29300
rect 11572 29288 11578 29300
rect 12621 29291 12679 29297
rect 12621 29288 12633 29291
rect 11572 29260 12633 29288
rect 11572 29248 11578 29260
rect 12621 29257 12633 29260
rect 12667 29257 12679 29291
rect 12621 29251 12679 29257
rect 15102 29248 15108 29300
rect 15160 29288 15166 29300
rect 15562 29288 15568 29300
rect 15160 29260 15568 29288
rect 15160 29248 15166 29260
rect 15562 29248 15568 29260
rect 15620 29248 15626 29300
rect 16850 29248 16856 29300
rect 16908 29288 16914 29300
rect 19981 29291 20039 29297
rect 19981 29288 19993 29291
rect 16908 29260 19993 29288
rect 16908 29248 16914 29260
rect 19981 29257 19993 29260
rect 20027 29257 20039 29291
rect 19981 29251 20039 29257
rect 20073 29291 20131 29297
rect 20073 29257 20085 29291
rect 20119 29288 20131 29291
rect 20530 29288 20536 29300
rect 20119 29260 20536 29288
rect 20119 29257 20131 29260
rect 20073 29251 20131 29257
rect 20530 29248 20536 29260
rect 20588 29248 20594 29300
rect 22462 29248 22468 29300
rect 22520 29248 22526 29300
rect 23661 29291 23719 29297
rect 23661 29257 23673 29291
rect 23707 29288 23719 29291
rect 24118 29288 24124 29300
rect 23707 29260 24124 29288
rect 23707 29257 23719 29260
rect 23661 29251 23719 29257
rect 24118 29248 24124 29260
rect 24176 29288 24182 29300
rect 25774 29288 25780 29300
rect 24176 29260 25780 29288
rect 24176 29248 24182 29260
rect 25774 29248 25780 29260
rect 25832 29248 25838 29300
rect 9677 29223 9735 29229
rect 9677 29189 9689 29223
rect 9723 29220 9735 29223
rect 9766 29220 9772 29232
rect 9723 29192 9772 29220
rect 9723 29189 9735 29192
rect 9677 29183 9735 29189
rect 9766 29180 9772 29192
rect 9824 29180 9830 29232
rect 11698 29220 11704 29232
rect 10902 29192 11704 29220
rect 11698 29180 11704 29192
rect 11756 29220 11762 29232
rect 13814 29220 13820 29232
rect 11756 29192 13820 29220
rect 11756 29180 11762 29192
rect 13814 29180 13820 29192
rect 13872 29180 13878 29232
rect 15841 29223 15899 29229
rect 15841 29189 15853 29223
rect 15887 29220 15899 29223
rect 15930 29220 15936 29232
rect 15887 29192 15936 29220
rect 15887 29189 15899 29192
rect 15841 29183 15899 29189
rect 15930 29180 15936 29192
rect 15988 29180 15994 29232
rect 17402 29180 17408 29232
rect 17460 29220 17466 29232
rect 21453 29223 21511 29229
rect 21453 29220 21465 29223
rect 17460 29192 21465 29220
rect 17460 29180 17466 29192
rect 21453 29189 21465 29192
rect 21499 29189 21511 29223
rect 21453 29183 21511 29189
rect 22373 29223 22431 29229
rect 22373 29189 22385 29223
rect 22419 29220 22431 29223
rect 24946 29220 24952 29232
rect 22419 29192 24952 29220
rect 22419 29189 22431 29192
rect 22373 29183 22431 29189
rect 24946 29180 24952 29192
rect 25004 29180 25010 29232
rect 11882 29112 11888 29164
rect 11940 29152 11946 29164
rect 11977 29155 12035 29161
rect 11977 29152 11989 29155
rect 11940 29124 11989 29152
rect 11940 29112 11946 29124
rect 11977 29121 11989 29124
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 12618 29112 12624 29164
rect 12676 29152 12682 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 12676 29124 13093 29152
rect 12676 29112 12682 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 16206 29112 16212 29164
rect 16264 29152 16270 29164
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 16264 29124 16865 29152
rect 16264 29112 16270 29124
rect 16853 29121 16865 29124
rect 16899 29121 16911 29155
rect 17945 29155 18003 29161
rect 17945 29152 17957 29155
rect 16853 29115 16911 29121
rect 17880 29124 17957 29152
rect 9398 29044 9404 29096
rect 9456 29044 9462 29096
rect 13998 29044 14004 29096
rect 14056 29084 14062 29096
rect 14829 29087 14887 29093
rect 14829 29084 14841 29087
rect 14056 29056 14841 29084
rect 14056 29044 14062 29056
rect 14829 29053 14841 29056
rect 14875 29053 14887 29087
rect 14829 29047 14887 29053
rect 15654 29044 15660 29096
rect 15712 29084 15718 29096
rect 15933 29087 15991 29093
rect 15933 29084 15945 29087
rect 15712 29056 15945 29084
rect 15712 29044 15718 29056
rect 15933 29053 15945 29056
rect 15979 29053 15991 29087
rect 15933 29047 15991 29053
rect 11146 28976 11152 29028
rect 11204 28976 11210 29028
rect 15948 29016 15976 29047
rect 16114 29044 16120 29096
rect 16172 29044 16178 29096
rect 16390 29044 16396 29096
rect 16448 29084 16454 29096
rect 16448 29056 17816 29084
rect 16448 29044 16454 29056
rect 16482 29016 16488 29028
rect 14752 28988 15608 29016
rect 15948 28988 16488 29016
rect 13344 28951 13402 28957
rect 13344 28917 13356 28951
rect 13390 28948 13402 28951
rect 14752 28948 14780 28988
rect 13390 28920 14780 28948
rect 13390 28917 13402 28920
rect 13344 28911 13402 28917
rect 15470 28908 15476 28960
rect 15528 28908 15534 28960
rect 15580 28948 15608 28988
rect 16482 28976 16488 28988
rect 16540 28976 16546 29028
rect 17788 28960 17816 29056
rect 17880 29016 17908 29124
rect 17945 29121 17957 29124
rect 17991 29121 18003 29155
rect 17945 29115 18003 29121
rect 18690 29112 18696 29164
rect 18748 29152 18754 29164
rect 20714 29152 20720 29164
rect 18748 29124 20720 29152
rect 18748 29112 18754 29124
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 20806 29112 20812 29164
rect 20864 29112 20870 29164
rect 22830 29112 22836 29164
rect 22888 29152 22894 29164
rect 22888 29124 23520 29152
rect 22888 29112 22894 29124
rect 19337 29087 19395 29093
rect 19337 29084 19349 29087
rect 18064 29056 19349 29084
rect 17954 29016 17960 29028
rect 17880 28988 17960 29016
rect 17954 28976 17960 28988
rect 18012 28976 18018 29028
rect 17497 28951 17555 28957
rect 17497 28948 17509 28951
rect 15580 28920 17509 28948
rect 17497 28917 17509 28920
rect 17543 28917 17555 28951
rect 17497 28911 17555 28917
rect 17770 28908 17776 28960
rect 17828 28948 17834 28960
rect 18064 28948 18092 29056
rect 19337 29053 19349 29056
rect 19383 29053 19395 29087
rect 19337 29047 19395 29053
rect 20257 29087 20315 29093
rect 20257 29053 20269 29087
rect 20303 29084 20315 29087
rect 21174 29084 21180 29096
rect 20303 29056 21180 29084
rect 20303 29053 20315 29056
rect 20257 29047 20315 29053
rect 21174 29044 21180 29056
rect 21232 29044 21238 29096
rect 22649 29087 22707 29093
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23382 29084 23388 29096
rect 22695 29056 23388 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23382 29044 23388 29056
rect 23440 29044 23446 29096
rect 23492 29084 23520 29124
rect 23566 29112 23572 29164
rect 23624 29152 23630 29164
rect 23624 29124 23888 29152
rect 23624 29112 23630 29124
rect 23753 29087 23811 29093
rect 23753 29084 23765 29087
rect 23492 29056 23765 29084
rect 23753 29053 23765 29056
rect 23799 29053 23811 29087
rect 23860 29084 23888 29124
rect 24394 29112 24400 29164
rect 24452 29112 24458 29164
rect 23934 29084 23940 29096
rect 23860 29056 23940 29084
rect 23753 29047 23811 29053
rect 23934 29044 23940 29056
rect 23992 29084 23998 29096
rect 24578 29084 24584 29096
rect 23992 29056 24584 29084
rect 23992 29044 23998 29056
rect 24578 29044 24584 29056
rect 24636 29044 24642 29096
rect 18230 28976 18236 29028
rect 18288 28976 18294 29028
rect 18322 28976 18328 29028
rect 18380 29016 18386 29028
rect 18601 29019 18659 29025
rect 18601 29016 18613 29019
rect 18380 28988 18613 29016
rect 18380 28976 18386 28988
rect 18601 28985 18613 28988
rect 18647 28985 18659 29019
rect 18601 28979 18659 28985
rect 18690 28976 18696 29028
rect 18748 29016 18754 29028
rect 19613 29019 19671 29025
rect 19613 29016 19625 29019
rect 18748 28988 19625 29016
rect 18748 28976 18754 28988
rect 19613 28985 19625 28988
rect 19659 28985 19671 29019
rect 19613 28979 19671 28985
rect 22002 28976 22008 29028
rect 22060 28976 22066 29028
rect 23198 28976 23204 29028
rect 23256 28976 23262 29028
rect 23290 28976 23296 29028
rect 23348 29016 23354 29028
rect 25041 29019 25099 29025
rect 25041 29016 25053 29019
rect 23348 28988 25053 29016
rect 23348 28976 23354 28988
rect 25041 28985 25053 28988
rect 25087 28985 25099 29019
rect 25041 28979 25099 28985
rect 17828 28920 18092 28948
rect 18248 28948 18276 28976
rect 18877 28951 18935 28957
rect 18877 28948 18889 28951
rect 18248 28920 18889 28948
rect 17828 28908 17834 28920
rect 18877 28917 18889 28920
rect 18923 28917 18935 28951
rect 18877 28911 18935 28917
rect 19153 28951 19211 28957
rect 19153 28917 19165 28951
rect 19199 28948 19211 28951
rect 19242 28948 19248 28960
rect 19199 28920 19248 28948
rect 19199 28917 19211 28920
rect 19153 28911 19211 28917
rect 19242 28908 19248 28920
rect 19300 28908 19306 28960
rect 19886 28908 19892 28960
rect 19944 28948 19950 28960
rect 22462 28948 22468 28960
rect 19944 28920 22468 28948
rect 19944 28908 19950 28920
rect 22462 28908 22468 28920
rect 22520 28908 22526 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 8846 28704 8852 28756
rect 8904 28744 8910 28756
rect 9677 28747 9735 28753
rect 9677 28744 9689 28747
rect 8904 28716 9689 28744
rect 8904 28704 8910 28716
rect 9677 28713 9689 28716
rect 9723 28713 9735 28747
rect 9677 28707 9735 28713
rect 12710 28704 12716 28756
rect 12768 28744 12774 28756
rect 12805 28747 12863 28753
rect 12805 28744 12817 28747
rect 12768 28716 12817 28744
rect 12768 28704 12774 28716
rect 12805 28713 12817 28716
rect 12851 28713 12863 28747
rect 14918 28744 14924 28756
rect 12805 28707 12863 28713
rect 13556 28716 14924 28744
rect 10686 28676 10692 28688
rect 7944 28648 10692 28676
rect 7944 28549 7972 28648
rect 10686 28636 10692 28648
rect 10744 28636 10750 28688
rect 10226 28568 10232 28620
rect 10284 28568 10290 28620
rect 11422 28568 11428 28620
rect 11480 28608 11486 28620
rect 13556 28617 13584 28716
rect 14918 28704 14924 28716
rect 14976 28704 14982 28756
rect 15304 28716 15608 28744
rect 15304 28676 15332 28716
rect 13648 28648 15332 28676
rect 15473 28679 15531 28685
rect 13541 28611 13599 28617
rect 11480 28580 13492 28608
rect 11480 28568 11486 28580
rect 7929 28543 7987 28549
rect 7929 28509 7941 28543
rect 7975 28509 7987 28543
rect 7929 28503 7987 28509
rect 8662 28500 8668 28552
rect 8720 28540 8726 28552
rect 9398 28540 9404 28552
rect 8720 28512 9404 28540
rect 8720 28500 8726 28512
rect 9398 28500 9404 28512
rect 9456 28540 9462 28552
rect 11054 28540 11060 28552
rect 9456 28512 11060 28540
rect 9456 28500 9462 28512
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 13464 28540 13492 28580
rect 13541 28577 13553 28611
rect 13587 28577 13599 28611
rect 13541 28571 13599 28577
rect 13648 28540 13676 28648
rect 15473 28645 15485 28679
rect 15519 28645 15531 28679
rect 15580 28676 15608 28716
rect 22370 28704 22376 28756
rect 22428 28744 22434 28756
rect 23845 28747 23903 28753
rect 22428 28716 23704 28744
rect 22428 28704 22434 28716
rect 17865 28679 17923 28685
rect 17865 28676 17877 28679
rect 15580 28648 17877 28676
rect 15473 28639 15531 28645
rect 17865 28645 17877 28648
rect 17911 28645 17923 28679
rect 23014 28676 23020 28688
rect 17865 28639 17923 28645
rect 17972 28648 23020 28676
rect 14734 28568 14740 28620
rect 14792 28568 14798 28620
rect 14829 28611 14887 28617
rect 14829 28577 14841 28611
rect 14875 28577 14887 28611
rect 14829 28571 14887 28577
rect 13464 28512 13676 28540
rect 13906 28500 13912 28552
rect 13964 28540 13970 28552
rect 14458 28540 14464 28552
rect 13964 28512 14464 28540
rect 13964 28500 13970 28512
rect 14458 28500 14464 28512
rect 14516 28540 14522 28552
rect 14844 28540 14872 28571
rect 15488 28540 15516 28639
rect 15930 28568 15936 28620
rect 15988 28568 15994 28620
rect 16022 28568 16028 28620
rect 16080 28568 16086 28620
rect 16850 28568 16856 28620
rect 16908 28608 16914 28620
rect 17221 28611 17279 28617
rect 17221 28608 17233 28611
rect 16908 28580 17233 28608
rect 16908 28568 16914 28580
rect 17221 28577 17233 28580
rect 17267 28577 17279 28611
rect 17221 28571 17279 28577
rect 17310 28568 17316 28620
rect 17368 28608 17374 28620
rect 17972 28608 18000 28648
rect 23014 28636 23020 28648
rect 23072 28636 23078 28688
rect 17368 28580 18000 28608
rect 18509 28611 18567 28617
rect 17368 28568 17374 28580
rect 18509 28577 18521 28611
rect 18555 28608 18567 28611
rect 18782 28608 18788 28620
rect 18555 28580 18788 28608
rect 18555 28577 18567 28580
rect 18509 28571 18567 28577
rect 18782 28568 18788 28580
rect 18840 28568 18846 28620
rect 21174 28568 21180 28620
rect 21232 28608 21238 28620
rect 22741 28611 22799 28617
rect 22741 28608 22753 28611
rect 21232 28580 22753 28608
rect 21232 28568 21238 28580
rect 22741 28577 22753 28580
rect 22787 28577 22799 28611
rect 23676 28608 23704 28716
rect 23845 28713 23857 28747
rect 23891 28744 23903 28747
rect 23934 28744 23940 28756
rect 23891 28716 23940 28744
rect 23891 28713 23903 28716
rect 23845 28707 23903 28713
rect 23934 28704 23940 28716
rect 23992 28704 23998 28756
rect 24118 28704 24124 28756
rect 24176 28704 24182 28756
rect 25041 28611 25099 28617
rect 25041 28608 25053 28611
rect 23676 28580 25053 28608
rect 22741 28571 22799 28577
rect 25041 28577 25053 28580
rect 25087 28577 25099 28611
rect 25041 28571 25099 28577
rect 25133 28611 25191 28617
rect 25133 28577 25145 28611
rect 25179 28577 25191 28611
rect 25133 28571 25191 28577
rect 14516 28512 14872 28540
rect 14936 28512 15516 28540
rect 15841 28543 15899 28549
rect 14516 28500 14522 28512
rect 8573 28475 8631 28481
rect 8573 28441 8585 28475
rect 8619 28472 8631 28475
rect 10502 28472 10508 28484
rect 8619 28444 10508 28472
rect 8619 28441 8631 28444
rect 8573 28435 8631 28441
rect 10502 28432 10508 28444
rect 10560 28432 10566 28484
rect 11330 28432 11336 28484
rect 11388 28432 11394 28484
rect 11790 28472 11796 28484
rect 11716 28444 11796 28472
rect 9950 28364 9956 28416
rect 10008 28404 10014 28416
rect 10045 28407 10103 28413
rect 10045 28404 10057 28407
rect 10008 28376 10057 28404
rect 10008 28364 10014 28376
rect 10045 28373 10057 28376
rect 10091 28373 10103 28407
rect 10045 28367 10103 28373
rect 10137 28407 10195 28413
rect 10137 28373 10149 28407
rect 10183 28404 10195 28407
rect 10410 28404 10416 28416
rect 10183 28376 10416 28404
rect 10183 28373 10195 28376
rect 10137 28367 10195 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 11716 28404 11744 28444
rect 11790 28432 11796 28444
rect 11848 28432 11854 28484
rect 13446 28432 13452 28484
rect 13504 28472 13510 28484
rect 14936 28472 14964 28512
rect 15841 28509 15853 28543
rect 15887 28509 15899 28543
rect 15841 28503 15899 28509
rect 13504 28444 14964 28472
rect 13504 28432 13510 28444
rect 15470 28432 15476 28484
rect 15528 28472 15534 28484
rect 15856 28472 15884 28503
rect 16666 28500 16672 28552
rect 16724 28540 16730 28552
rect 17037 28543 17095 28549
rect 16724 28512 16804 28540
rect 16724 28500 16730 28512
rect 15528 28444 15884 28472
rect 15528 28432 15534 28444
rect 13173 28407 13231 28413
rect 13173 28404 13185 28407
rect 11716 28376 13185 28404
rect 13173 28373 13185 28376
rect 13219 28373 13231 28407
rect 13173 28367 13231 28373
rect 13630 28364 13636 28416
rect 13688 28404 13694 28416
rect 14277 28407 14335 28413
rect 14277 28404 14289 28407
rect 13688 28376 14289 28404
rect 13688 28364 13694 28376
rect 14277 28373 14289 28376
rect 14323 28373 14335 28407
rect 14277 28367 14335 28373
rect 14645 28407 14703 28413
rect 14645 28373 14657 28407
rect 14691 28404 14703 28407
rect 16574 28404 16580 28416
rect 14691 28376 16580 28404
rect 14691 28373 14703 28376
rect 14645 28367 14703 28373
rect 16574 28364 16580 28376
rect 16632 28364 16638 28416
rect 16666 28364 16672 28416
rect 16724 28364 16730 28416
rect 16776 28404 16804 28512
rect 17037 28509 17049 28543
rect 17083 28540 17095 28543
rect 17770 28540 17776 28552
rect 17083 28512 17776 28540
rect 17083 28509 17095 28512
rect 17037 28503 17095 28509
rect 17770 28500 17776 28512
rect 17828 28500 17834 28552
rect 18325 28543 18383 28549
rect 18325 28509 18337 28543
rect 18371 28540 18383 28543
rect 19518 28540 19524 28552
rect 18371 28512 19524 28540
rect 18371 28509 18383 28512
rect 18325 28503 18383 28509
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 20809 28543 20867 28549
rect 20809 28509 20821 28543
rect 20855 28540 20867 28543
rect 20855 28512 21956 28540
rect 20855 28509 20867 28512
rect 20809 28503 20867 28509
rect 21928 28484 21956 28512
rect 22462 28500 22468 28552
rect 22520 28540 22526 28552
rect 22649 28543 22707 28549
rect 22649 28540 22661 28543
rect 22520 28512 22661 28540
rect 22520 28500 22526 28512
rect 22649 28509 22661 28512
rect 22695 28509 22707 28543
rect 22649 28503 22707 28509
rect 23566 28500 23572 28552
rect 23624 28540 23630 28552
rect 25148 28540 25176 28571
rect 23624 28512 25176 28540
rect 23624 28500 23630 28512
rect 16942 28432 16948 28484
rect 17000 28472 17006 28484
rect 18233 28475 18291 28481
rect 18233 28472 18245 28475
rect 17000 28444 18245 28472
rect 17000 28432 17006 28444
rect 18233 28441 18245 28444
rect 18279 28441 18291 28475
rect 18233 28435 18291 28441
rect 18598 28432 18604 28484
rect 18656 28472 18662 28484
rect 19429 28475 19487 28481
rect 19429 28472 19441 28475
rect 18656 28444 19441 28472
rect 18656 28432 18662 28444
rect 19429 28441 19441 28444
rect 19475 28441 19487 28475
rect 19429 28435 19487 28441
rect 20162 28432 20168 28484
rect 20220 28432 20226 28484
rect 20438 28432 20444 28484
rect 20496 28472 20502 28484
rect 21545 28475 21603 28481
rect 21545 28472 21557 28475
rect 20496 28444 21557 28472
rect 20496 28432 20502 28444
rect 21545 28441 21557 28444
rect 21591 28441 21603 28475
rect 21545 28435 21603 28441
rect 21910 28432 21916 28484
rect 21968 28472 21974 28484
rect 23201 28475 23259 28481
rect 23201 28472 23213 28475
rect 21968 28444 23213 28472
rect 21968 28432 21974 28444
rect 23201 28441 23213 28444
rect 23247 28472 23259 28475
rect 23385 28475 23443 28481
rect 23385 28472 23397 28475
rect 23247 28444 23397 28472
rect 23247 28441 23259 28444
rect 23201 28435 23259 28441
rect 23385 28441 23397 28444
rect 23431 28441 23443 28475
rect 23385 28435 23443 28441
rect 23661 28475 23719 28481
rect 23661 28441 23673 28475
rect 23707 28472 23719 28475
rect 24394 28472 24400 28484
rect 23707 28444 24400 28472
rect 23707 28441 23719 28444
rect 23661 28435 23719 28441
rect 17129 28407 17187 28413
rect 17129 28404 17141 28407
rect 16776 28376 17141 28404
rect 17129 28373 17141 28376
rect 17175 28404 17187 28407
rect 17310 28404 17316 28416
rect 17175 28376 17316 28404
rect 17175 28373 17187 28376
rect 17129 28367 17187 28373
rect 17310 28364 17316 28376
rect 17368 28404 17374 28416
rect 18877 28407 18935 28413
rect 18877 28404 18889 28407
rect 17368 28376 18889 28404
rect 17368 28364 17374 28376
rect 18877 28373 18889 28376
rect 18923 28373 18935 28407
rect 18877 28367 18935 28373
rect 22186 28364 22192 28416
rect 22244 28364 22250 28416
rect 22557 28407 22615 28413
rect 22557 28373 22569 28407
rect 22603 28404 22615 28407
rect 23676 28404 23704 28435
rect 24394 28432 24400 28444
rect 24452 28472 24458 28484
rect 25774 28472 25780 28484
rect 24452 28444 25780 28472
rect 24452 28432 24458 28444
rect 25774 28432 25780 28444
rect 25832 28432 25838 28484
rect 22603 28376 23704 28404
rect 22603 28373 22615 28376
rect 22557 28367 22615 28373
rect 23750 28364 23756 28416
rect 23808 28404 23814 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 23808 28376 24593 28404
rect 23808 28364 23814 28376
rect 24581 28373 24593 28376
rect 24627 28373 24639 28407
rect 24581 28367 24639 28373
rect 24762 28364 24768 28416
rect 24820 28404 24826 28416
rect 24949 28407 25007 28413
rect 24949 28404 24961 28407
rect 24820 28376 24961 28404
rect 24820 28364 24826 28376
rect 24949 28373 24961 28376
rect 24995 28373 25007 28407
rect 24949 28367 25007 28373
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 10226 28160 10232 28212
rect 10284 28200 10290 28212
rect 10413 28203 10471 28209
rect 10413 28200 10425 28203
rect 10284 28172 10425 28200
rect 10284 28160 10290 28172
rect 10413 28169 10425 28172
rect 10459 28169 10471 28203
rect 10413 28163 10471 28169
rect 10689 28203 10747 28209
rect 10689 28169 10701 28203
rect 10735 28200 10747 28203
rect 11241 28203 11299 28209
rect 11241 28200 11253 28203
rect 10735 28172 11253 28200
rect 10735 28169 10747 28172
rect 10689 28163 10747 28169
rect 11241 28169 11253 28172
rect 11287 28200 11299 28203
rect 11698 28200 11704 28212
rect 11287 28172 11704 28200
rect 11287 28169 11299 28172
rect 11241 28163 11299 28169
rect 10704 28132 10732 28163
rect 11698 28160 11704 28172
rect 11756 28160 11762 28212
rect 13541 28203 13599 28209
rect 13541 28169 13553 28203
rect 13587 28200 13599 28203
rect 14642 28200 14648 28212
rect 13587 28172 14648 28200
rect 13587 28169 13599 28172
rect 13541 28163 13599 28169
rect 14642 28160 14648 28172
rect 14700 28200 14706 28212
rect 15749 28203 15807 28209
rect 14700 28172 15608 28200
rect 14700 28160 14706 28172
rect 10166 28104 10732 28132
rect 11716 28132 11744 28160
rect 14366 28132 14372 28144
rect 11716 28104 12558 28132
rect 14016 28104 14372 28132
rect 8662 28024 8668 28076
rect 8720 28024 8726 28076
rect 11054 28024 11060 28076
rect 11112 28064 11118 28076
rect 14016 28073 14044 28104
rect 14366 28092 14372 28104
rect 14424 28092 14430 28144
rect 15286 28092 15292 28144
rect 15344 28092 15350 28144
rect 15580 28132 15608 28172
rect 15749 28169 15761 28203
rect 15795 28200 15807 28203
rect 16850 28200 16856 28212
rect 15795 28172 16856 28200
rect 15795 28169 15807 28172
rect 15749 28163 15807 28169
rect 16850 28160 16856 28172
rect 16908 28160 16914 28212
rect 16942 28160 16948 28212
rect 17000 28160 17006 28212
rect 19334 28160 19340 28212
rect 19392 28160 19398 28212
rect 20441 28203 20499 28209
rect 20441 28169 20453 28203
rect 20487 28200 20499 28203
rect 20806 28200 20812 28212
rect 20487 28172 20812 28200
rect 20487 28169 20499 28172
rect 20441 28163 20499 28169
rect 20806 28160 20812 28172
rect 20864 28160 20870 28212
rect 24949 28203 25007 28209
rect 24949 28169 24961 28203
rect 24995 28200 25007 28203
rect 25038 28200 25044 28212
rect 24995 28172 25044 28200
rect 24995 28169 25007 28172
rect 24949 28163 25007 28169
rect 25038 28160 25044 28172
rect 25096 28160 25102 28212
rect 17862 28132 17868 28144
rect 15580 28104 17868 28132
rect 17862 28092 17868 28104
rect 17920 28092 17926 28144
rect 18414 28092 18420 28144
rect 18472 28092 18478 28144
rect 22278 28092 22284 28144
rect 22336 28132 22342 28144
rect 22336 28104 22770 28132
rect 22336 28092 22342 28104
rect 11793 28067 11851 28073
rect 11793 28064 11805 28067
rect 11112 28036 11805 28064
rect 11112 28024 11118 28036
rect 11793 28033 11805 28036
rect 11839 28033 11851 28067
rect 11793 28027 11851 28033
rect 14001 28067 14059 28073
rect 14001 28033 14013 28067
rect 14047 28033 14059 28067
rect 14001 28027 14059 28033
rect 8938 27956 8944 28008
rect 8996 27956 9002 28008
rect 11808 27860 11836 28027
rect 12069 27999 12127 28005
rect 12069 27965 12081 27999
rect 12115 27996 12127 27999
rect 12434 27996 12440 28008
rect 12115 27968 12440 27996
rect 12115 27965 12127 27968
rect 12069 27959 12127 27965
rect 12434 27956 12440 27968
rect 12492 27956 12498 28008
rect 14016 27928 14044 28027
rect 17034 28024 17040 28076
rect 17092 28064 17098 28076
rect 17589 28067 17647 28073
rect 17589 28064 17601 28067
rect 17092 28036 17601 28064
rect 17092 28024 17098 28036
rect 17589 28033 17601 28036
rect 17635 28033 17647 28067
rect 17589 28027 17647 28033
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28064 19855 28067
rect 20898 28064 20904 28076
rect 19843 28036 20904 28064
rect 19843 28033 19855 28036
rect 19797 28027 19855 28033
rect 20898 28024 20904 28036
rect 20956 28024 20962 28076
rect 20993 28067 21051 28073
rect 20993 28033 21005 28067
rect 21039 28064 21051 28067
rect 21266 28064 21272 28076
rect 21039 28036 21272 28064
rect 21039 28033 21051 28036
rect 20993 28027 21051 28033
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 22002 28024 22008 28076
rect 22060 28024 22066 28076
rect 24210 28024 24216 28076
rect 24268 28064 24274 28076
rect 25041 28067 25099 28073
rect 25041 28064 25053 28067
rect 24268 28036 25053 28064
rect 24268 28024 24274 28036
rect 25041 28033 25053 28036
rect 25087 28033 25099 28067
rect 25041 28027 25099 28033
rect 14277 27999 14335 28005
rect 14277 27996 14289 27999
rect 13464 27900 14044 27928
rect 14108 27968 14289 27996
rect 13464 27860 13492 27900
rect 11808 27832 13492 27860
rect 13722 27820 13728 27872
rect 13780 27860 13786 27872
rect 14108 27860 14136 27968
rect 14277 27965 14289 27968
rect 14323 27965 14335 27999
rect 14277 27959 14335 27965
rect 14918 27956 14924 28008
rect 14976 27996 14982 28008
rect 17865 27999 17923 28005
rect 14976 27968 17724 27996
rect 14976 27956 14982 27968
rect 13780 27832 14136 27860
rect 13780 27820 13786 27832
rect 15470 27820 15476 27872
rect 15528 27860 15534 27872
rect 15746 27860 15752 27872
rect 15528 27832 15752 27860
rect 15528 27820 15534 27832
rect 15746 27820 15752 27832
rect 15804 27860 15810 27872
rect 16114 27860 16120 27872
rect 15804 27832 16120 27860
rect 15804 27820 15810 27832
rect 16114 27820 16120 27832
rect 16172 27820 16178 27872
rect 16393 27863 16451 27869
rect 16393 27829 16405 27863
rect 16439 27860 16451 27863
rect 16482 27860 16488 27872
rect 16439 27832 16488 27860
rect 16439 27829 16451 27832
rect 16393 27823 16451 27829
rect 16482 27820 16488 27832
rect 16540 27820 16546 27872
rect 17696 27860 17724 27968
rect 17865 27965 17877 27999
rect 17911 27996 17923 27999
rect 20070 27996 20076 28008
rect 17911 27968 20076 27996
rect 17911 27965 17923 27968
rect 17865 27959 17923 27965
rect 20070 27956 20076 27968
rect 20128 27956 20134 28008
rect 21082 27956 21088 28008
rect 21140 27996 21146 28008
rect 21177 27999 21235 28005
rect 21177 27996 21189 27999
rect 21140 27968 21189 27996
rect 21140 27956 21146 27968
rect 21177 27965 21189 27968
rect 21223 27965 21235 27999
rect 21177 27959 21235 27965
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 22738 27996 22744 28008
rect 22327 27968 22744 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 22738 27956 22744 27968
rect 22796 27956 22802 28008
rect 25130 27956 25136 28008
rect 25188 27956 25194 28008
rect 19242 27888 19248 27940
rect 19300 27928 19306 27940
rect 21100 27928 21128 27956
rect 19300 27900 21128 27928
rect 19300 27888 19306 27900
rect 24578 27888 24584 27940
rect 24636 27888 24642 27940
rect 21910 27860 21916 27872
rect 17696 27832 21916 27860
rect 21910 27820 21916 27832
rect 21968 27820 21974 27872
rect 23014 27820 23020 27872
rect 23072 27860 23078 27872
rect 23382 27860 23388 27872
rect 23072 27832 23388 27860
rect 23072 27820 23078 27832
rect 23382 27820 23388 27832
rect 23440 27820 23446 27872
rect 23566 27820 23572 27872
rect 23624 27860 23630 27872
rect 23753 27863 23811 27869
rect 23753 27860 23765 27863
rect 23624 27832 23765 27860
rect 23624 27820 23630 27832
rect 23753 27829 23765 27832
rect 23799 27829 23811 27863
rect 23753 27823 23811 27829
rect 24026 27820 24032 27872
rect 24084 27860 24090 27872
rect 24121 27863 24179 27869
rect 24121 27860 24133 27863
rect 24084 27832 24133 27860
rect 24084 27820 24090 27832
rect 24121 27829 24133 27832
rect 24167 27860 24179 27863
rect 24762 27860 24768 27872
rect 24167 27832 24768 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 10124 27659 10182 27665
rect 10124 27625 10136 27659
rect 10170 27656 10182 27659
rect 10318 27656 10324 27668
rect 10170 27628 10324 27656
rect 10170 27625 10182 27628
rect 10124 27619 10182 27625
rect 10318 27616 10324 27628
rect 10376 27616 10382 27668
rect 11698 27616 11704 27668
rect 11756 27656 11762 27668
rect 11885 27659 11943 27665
rect 11885 27656 11897 27659
rect 11756 27628 11897 27656
rect 11756 27616 11762 27628
rect 11885 27625 11897 27628
rect 11931 27656 11943 27659
rect 14553 27659 14611 27665
rect 11931 27628 13860 27656
rect 11931 27625 11943 27628
rect 11885 27619 11943 27625
rect 13722 27548 13728 27600
rect 13780 27548 13786 27600
rect 13832 27588 13860 27628
rect 14553 27625 14565 27659
rect 14599 27656 14611 27659
rect 16482 27656 16488 27668
rect 14599 27628 16488 27656
rect 14599 27625 14611 27628
rect 14553 27619 14611 27625
rect 16482 27616 16488 27628
rect 16540 27616 16546 27668
rect 18598 27616 18604 27668
rect 18656 27656 18662 27668
rect 20888 27659 20946 27665
rect 18656 27628 19656 27656
rect 18656 27616 18662 27628
rect 14185 27591 14243 27597
rect 14185 27588 14197 27591
rect 13832 27560 14197 27588
rect 14185 27557 14197 27560
rect 14231 27588 14243 27591
rect 15286 27588 15292 27600
rect 14231 27560 15292 27588
rect 14231 27557 14243 27560
rect 14185 27551 14243 27557
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 15396 27560 19564 27588
rect 9861 27523 9919 27529
rect 9861 27489 9873 27523
rect 9907 27520 9919 27523
rect 10870 27520 10876 27532
rect 9907 27492 10876 27520
rect 9907 27489 9919 27492
rect 9861 27483 9919 27489
rect 10870 27480 10876 27492
rect 10928 27480 10934 27532
rect 15396 27520 15424 27560
rect 12406 27492 15424 27520
rect 15473 27523 15531 27529
rect 11698 27384 11704 27396
rect 11362 27356 11704 27384
rect 11698 27344 11704 27356
rect 11756 27344 11762 27396
rect 12161 27387 12219 27393
rect 12161 27353 12173 27387
rect 12207 27384 12219 27387
rect 12406 27384 12434 27492
rect 12636 27461 12664 27492
rect 15473 27489 15485 27523
rect 15519 27489 15531 27523
rect 15473 27483 15531 27489
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27452 12679 27455
rect 13081 27455 13139 27461
rect 12667 27424 12701 27452
rect 12667 27421 12679 27424
rect 12621 27415 12679 27421
rect 13081 27421 13093 27455
rect 13127 27452 13139 27455
rect 15102 27452 15108 27464
rect 13127 27424 15108 27452
rect 13127 27421 13139 27424
rect 13081 27415 13139 27421
rect 15102 27412 15108 27424
rect 15160 27412 15166 27464
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27452 15255 27455
rect 15286 27452 15292 27464
rect 15243 27424 15292 27452
rect 15243 27421 15255 27424
rect 15197 27415 15255 27421
rect 15286 27412 15292 27424
rect 15344 27412 15350 27464
rect 15488 27452 15516 27483
rect 15930 27480 15936 27532
rect 15988 27520 15994 27532
rect 16577 27523 16635 27529
rect 16577 27520 16589 27523
rect 15988 27492 16589 27520
rect 15988 27480 15994 27492
rect 16577 27489 16589 27492
rect 16623 27489 16635 27523
rect 16577 27483 16635 27489
rect 16850 27480 16856 27532
rect 16908 27520 16914 27532
rect 17773 27523 17831 27529
rect 17773 27520 17785 27523
rect 16908 27492 17785 27520
rect 16908 27480 16914 27492
rect 17773 27489 17785 27492
rect 17819 27489 17831 27523
rect 19242 27520 19248 27532
rect 17773 27483 17831 27489
rect 18524 27492 19248 27520
rect 16758 27452 16764 27464
rect 15396 27424 15516 27452
rect 15672 27424 16764 27452
rect 12207 27356 12434 27384
rect 12207 27353 12219 27356
rect 12161 27347 12219 27353
rect 13998 27344 14004 27396
rect 14056 27384 14062 27396
rect 15396 27384 15424 27424
rect 14056 27356 15424 27384
rect 14056 27344 14062 27356
rect 9125 27319 9183 27325
rect 9125 27285 9137 27319
rect 9171 27316 9183 27319
rect 9306 27316 9312 27328
rect 9171 27288 9312 27316
rect 9171 27285 9183 27288
rect 9125 27279 9183 27285
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 11606 27276 11612 27328
rect 11664 27276 11670 27328
rect 12437 27319 12495 27325
rect 12437 27285 12449 27319
rect 12483 27316 12495 27319
rect 13722 27316 13728 27328
rect 12483 27288 13728 27316
rect 12483 27285 12495 27288
rect 12437 27279 12495 27285
rect 13722 27276 13728 27288
rect 13780 27276 13786 27328
rect 14369 27319 14427 27325
rect 14369 27285 14381 27319
rect 14415 27316 14427 27319
rect 14734 27316 14740 27328
rect 14415 27288 14740 27316
rect 14415 27285 14427 27288
rect 14369 27279 14427 27285
rect 14734 27276 14740 27288
rect 14792 27276 14798 27328
rect 14826 27276 14832 27328
rect 14884 27276 14890 27328
rect 15289 27319 15347 27325
rect 15289 27285 15301 27319
rect 15335 27316 15347 27319
rect 15672 27316 15700 27424
rect 16758 27412 16764 27424
rect 16816 27412 16822 27464
rect 17586 27412 17592 27464
rect 17644 27412 17650 27464
rect 18524 27461 18552 27492
rect 19242 27480 19248 27492
rect 19300 27480 19306 27532
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27421 18567 27455
rect 18509 27415 18567 27421
rect 15746 27344 15752 27396
rect 15804 27384 15810 27396
rect 15804 27356 16068 27384
rect 15804 27344 15810 27356
rect 16040 27325 16068 27356
rect 16206 27344 16212 27396
rect 16264 27384 16270 27396
rect 18524 27384 18552 27415
rect 18598 27412 18604 27464
rect 18656 27452 18662 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 18656 27424 19441 27452
rect 18656 27412 18662 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 16264 27356 18552 27384
rect 16264 27344 16270 27356
rect 15335 27288 15700 27316
rect 16025 27319 16083 27325
rect 15335 27285 15347 27288
rect 15289 27279 15347 27285
rect 16025 27285 16037 27319
rect 16071 27285 16083 27319
rect 16025 27279 16083 27285
rect 16298 27276 16304 27328
rect 16356 27316 16362 27328
rect 16393 27319 16451 27325
rect 16393 27316 16405 27319
rect 16356 27288 16405 27316
rect 16356 27276 16362 27288
rect 16393 27285 16405 27288
rect 16439 27285 16451 27319
rect 16393 27279 16451 27285
rect 16482 27276 16488 27328
rect 16540 27276 16546 27328
rect 16574 27276 16580 27328
rect 16632 27316 16638 27328
rect 17221 27319 17279 27325
rect 17221 27316 17233 27319
rect 16632 27288 17233 27316
rect 16632 27276 16638 27288
rect 17221 27285 17233 27288
rect 17267 27285 17279 27319
rect 17221 27279 17279 27285
rect 17681 27319 17739 27325
rect 17681 27285 17693 27319
rect 17727 27316 17739 27319
rect 18782 27316 18788 27328
rect 17727 27288 18788 27316
rect 17727 27285 17739 27288
rect 17681 27279 17739 27285
rect 18782 27276 18788 27288
rect 18840 27276 18846 27328
rect 19536 27316 19564 27560
rect 19628 27384 19656 27628
rect 20888 27625 20900 27659
rect 20934 27656 20946 27659
rect 23290 27656 23296 27668
rect 20934 27628 23296 27656
rect 20934 27625 20946 27628
rect 20888 27619 20946 27625
rect 23290 27616 23296 27628
rect 23348 27616 23354 27668
rect 23474 27616 23480 27668
rect 23532 27656 23538 27668
rect 23750 27656 23756 27668
rect 23532 27628 23756 27656
rect 23532 27616 23538 27628
rect 23750 27616 23756 27628
rect 23808 27616 23814 27668
rect 20070 27548 20076 27600
rect 20128 27548 20134 27600
rect 21910 27548 21916 27600
rect 21968 27588 21974 27600
rect 21968 27560 23244 27588
rect 21968 27548 21974 27560
rect 19702 27480 19708 27532
rect 19760 27520 19766 27532
rect 19760 27492 23152 27520
rect 19760 27480 19766 27492
rect 20438 27412 20444 27464
rect 20496 27452 20502 27464
rect 20625 27455 20683 27461
rect 20625 27452 20637 27455
rect 20496 27424 20637 27452
rect 20496 27412 20502 27424
rect 20625 27421 20637 27424
rect 20671 27421 20683 27455
rect 20625 27415 20683 27421
rect 22922 27384 22928 27396
rect 19628 27356 21390 27384
rect 22388 27356 22928 27384
rect 22278 27316 22284 27328
rect 19536 27288 22284 27316
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 22388 27325 22416 27356
rect 22922 27344 22928 27356
rect 22980 27344 22986 27396
rect 23124 27384 23152 27492
rect 23216 27461 23244 27560
rect 24872 27560 25176 27588
rect 23385 27523 23443 27529
rect 23385 27489 23397 27523
rect 23431 27520 23443 27523
rect 24486 27520 24492 27532
rect 23431 27492 24492 27520
rect 23431 27489 23443 27492
rect 23385 27483 23443 27489
rect 24486 27480 24492 27492
rect 24544 27480 24550 27532
rect 24872 27520 24900 27560
rect 25148 27529 25176 27560
rect 24780 27492 24900 27520
rect 25133 27523 25191 27529
rect 23201 27455 23259 27461
rect 23201 27421 23213 27455
rect 23247 27421 23259 27455
rect 23201 27415 23259 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27452 23351 27455
rect 23842 27452 23848 27464
rect 23339 27424 23848 27452
rect 23339 27421 23351 27424
rect 23293 27415 23351 27421
rect 23842 27412 23848 27424
rect 23900 27412 23906 27464
rect 24302 27412 24308 27464
rect 24360 27452 24366 27464
rect 24780 27452 24808 27492
rect 25133 27489 25145 27523
rect 25179 27489 25191 27523
rect 25133 27483 25191 27489
rect 24360 27424 24808 27452
rect 24360 27412 24366 27424
rect 25041 27387 25099 27393
rect 25041 27384 25053 27387
rect 23124 27356 25053 27384
rect 25041 27353 25053 27356
rect 25087 27353 25099 27387
rect 25041 27347 25099 27353
rect 22373 27319 22431 27325
rect 22373 27285 22385 27319
rect 22419 27285 22431 27319
rect 22373 27279 22431 27285
rect 22830 27276 22836 27328
rect 22888 27276 22894 27328
rect 24118 27276 24124 27328
rect 24176 27276 24182 27328
rect 24210 27276 24216 27328
rect 24268 27316 24274 27328
rect 24581 27319 24639 27325
rect 24581 27316 24593 27319
rect 24268 27288 24593 27316
rect 24268 27276 24274 27288
rect 24581 27285 24593 27288
rect 24627 27285 24639 27319
rect 24581 27279 24639 27285
rect 24946 27276 24952 27328
rect 25004 27276 25010 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 11149 27115 11207 27121
rect 11149 27081 11161 27115
rect 11195 27112 11207 27115
rect 11330 27112 11336 27124
rect 11195 27084 11336 27112
rect 11195 27081 11207 27084
rect 11149 27075 11207 27081
rect 11330 27072 11336 27084
rect 11388 27072 11394 27124
rect 12434 27072 12440 27124
rect 12492 27112 12498 27124
rect 12529 27115 12587 27121
rect 12529 27112 12541 27115
rect 12492 27084 12541 27112
rect 12492 27072 12498 27084
rect 12529 27081 12541 27084
rect 12575 27081 12587 27115
rect 12529 27075 12587 27081
rect 12989 27115 13047 27121
rect 12989 27081 13001 27115
rect 13035 27112 13047 27115
rect 13035 27084 16344 27112
rect 13035 27081 13047 27084
rect 12989 27075 13047 27081
rect 10226 27004 10232 27056
rect 10284 27044 10290 27056
rect 13357 27047 13415 27053
rect 13357 27044 13369 27047
rect 10284 27016 13369 27044
rect 10284 27004 10290 27016
rect 13357 27013 13369 27016
rect 13403 27013 13415 27047
rect 13357 27007 13415 27013
rect 13446 27004 13452 27056
rect 13504 27004 13510 27056
rect 13906 27004 13912 27056
rect 13964 27044 13970 27056
rect 15746 27044 15752 27056
rect 13964 27016 15752 27044
rect 13964 27004 13970 27016
rect 15746 27004 15752 27016
rect 15804 27004 15810 27056
rect 15841 27047 15899 27053
rect 15841 27013 15853 27047
rect 15887 27044 15899 27047
rect 16206 27044 16212 27056
rect 15887 27016 16212 27044
rect 15887 27013 15899 27016
rect 15841 27007 15899 27013
rect 8297 26979 8355 26985
rect 8297 26945 8309 26979
rect 8343 26976 8355 26979
rect 9306 26976 9312 26988
rect 8343 26948 9312 26976
rect 8343 26945 8355 26948
rect 8297 26939 8355 26945
rect 9306 26936 9312 26948
rect 9364 26936 9370 26988
rect 9398 26936 9404 26988
rect 9456 26936 9462 26988
rect 10502 26936 10508 26988
rect 10560 26936 10566 26988
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12066 26976 12072 26988
rect 11931 26948 12072 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12066 26936 12072 26948
rect 12124 26936 12130 26988
rect 15010 26976 15016 26988
rect 12406 26948 13584 26976
rect 4246 26868 4252 26920
rect 4304 26908 4310 26920
rect 10962 26908 10968 26920
rect 4304 26880 10968 26908
rect 4304 26868 4310 26880
rect 10962 26868 10968 26880
rect 11020 26868 11026 26920
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 12406 26908 12434 26948
rect 13556 26917 13584 26948
rect 14844 26948 15016 26976
rect 11204 26880 12434 26908
rect 13541 26911 13599 26917
rect 11204 26868 11210 26880
rect 13541 26877 13553 26911
rect 13587 26877 13599 26911
rect 13541 26871 13599 26877
rect 13354 26800 13360 26852
rect 13412 26840 13418 26852
rect 14737 26843 14795 26849
rect 14737 26840 14749 26843
rect 13412 26812 14749 26840
rect 13412 26800 13418 26812
rect 14737 26809 14749 26812
rect 14783 26809 14795 26843
rect 14737 26803 14795 26809
rect 6822 26732 6828 26784
rect 6880 26772 6886 26784
rect 8941 26775 8999 26781
rect 8941 26772 8953 26775
rect 6880 26744 8953 26772
rect 6880 26732 6886 26744
rect 8941 26741 8953 26744
rect 8987 26741 8999 26775
rect 8941 26735 8999 26741
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 10045 26775 10103 26781
rect 10045 26772 10057 26775
rect 9732 26744 10057 26772
rect 9732 26732 9738 26744
rect 10045 26741 10057 26744
rect 10091 26741 10103 26775
rect 10045 26735 10103 26741
rect 12250 26732 12256 26784
rect 12308 26772 12314 26784
rect 13998 26772 14004 26784
rect 12308 26744 14004 26772
rect 12308 26732 12314 26744
rect 13998 26732 14004 26744
rect 14056 26732 14062 26784
rect 14274 26732 14280 26784
rect 14332 26772 14338 26784
rect 14369 26775 14427 26781
rect 14369 26772 14381 26775
rect 14332 26744 14381 26772
rect 14332 26732 14338 26744
rect 14369 26741 14381 26744
rect 14415 26772 14427 26775
rect 14844 26772 14872 26948
rect 15010 26936 15016 26948
rect 15068 26976 15074 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 15068 26948 15117 26976
rect 15068 26936 15074 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 15197 26979 15255 26985
rect 15197 26945 15209 26979
rect 15243 26976 15255 26979
rect 15470 26976 15476 26988
rect 15243 26948 15476 26976
rect 15243 26945 15255 26948
rect 15197 26939 15255 26945
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 15562 26936 15568 26988
rect 15620 26976 15626 26988
rect 15856 26976 15884 27007
rect 16206 27004 16212 27016
rect 16264 27004 16270 27056
rect 16316 26985 16344 27084
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 19392 27084 20300 27112
rect 19392 27072 19398 27084
rect 16482 27004 16488 27056
rect 16540 27044 16546 27056
rect 17402 27044 17408 27056
rect 16540 27016 17408 27044
rect 16540 27004 16546 27016
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 20162 27044 20168 27056
rect 19550 27016 20168 27044
rect 20162 27004 20168 27016
rect 20220 27004 20226 27056
rect 15620 26948 15884 26976
rect 16301 26979 16359 26985
rect 15620 26936 15626 26948
rect 16301 26945 16313 26979
rect 16347 26945 16359 26979
rect 16301 26939 16359 26945
rect 16850 26936 16856 26988
rect 16908 26936 16914 26988
rect 17126 26936 17132 26988
rect 17184 26976 17190 26988
rect 17862 26976 17868 26988
rect 17184 26948 17868 26976
rect 17184 26936 17190 26948
rect 17862 26936 17868 26948
rect 17920 26976 17926 26988
rect 20272 26985 20300 27084
rect 20898 27072 20904 27124
rect 20956 27072 20962 27124
rect 21082 27072 21088 27124
rect 21140 27112 21146 27124
rect 21177 27115 21235 27121
rect 21177 27112 21189 27115
rect 21140 27084 21189 27112
rect 21140 27072 21146 27084
rect 21177 27081 21189 27084
rect 21223 27081 21235 27115
rect 21177 27075 21235 27081
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 21545 27115 21603 27121
rect 21545 27112 21557 27115
rect 21324 27084 21557 27112
rect 21324 27072 21330 27084
rect 21545 27081 21557 27084
rect 21591 27112 21603 27115
rect 21818 27112 21824 27124
rect 21591 27084 21824 27112
rect 21591 27081 21603 27084
rect 21545 27075 21603 27081
rect 21818 27072 21824 27084
rect 21876 27072 21882 27124
rect 22094 27072 22100 27124
rect 22152 27112 22158 27124
rect 22462 27112 22468 27124
rect 22152 27084 22468 27112
rect 22152 27072 22158 27084
rect 22462 27072 22468 27084
rect 22520 27112 22526 27124
rect 22520 27084 23428 27112
rect 22520 27072 22526 27084
rect 22370 27044 22376 27056
rect 21376 27016 22376 27044
rect 18049 26979 18107 26985
rect 18049 26976 18061 26979
rect 17920 26948 18061 26976
rect 17920 26936 17926 26948
rect 18049 26945 18061 26948
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 20257 26979 20315 26985
rect 20257 26945 20269 26979
rect 20303 26945 20315 26979
rect 20257 26939 20315 26945
rect 14918 26868 14924 26920
rect 14976 26908 14982 26920
rect 15381 26911 15439 26917
rect 15381 26908 15393 26911
rect 14976 26880 15393 26908
rect 14976 26868 14982 26880
rect 15381 26877 15393 26880
rect 15427 26908 15439 26911
rect 15930 26908 15936 26920
rect 15427 26880 15936 26908
rect 15427 26877 15439 26880
rect 15381 26871 15439 26877
rect 15930 26868 15936 26880
rect 15988 26868 15994 26920
rect 18325 26911 18383 26917
rect 18325 26877 18337 26911
rect 18371 26908 18383 26911
rect 21266 26908 21272 26920
rect 18371 26880 21272 26908
rect 18371 26877 18383 26880
rect 18325 26871 18383 26877
rect 21266 26868 21272 26880
rect 21324 26868 21330 26920
rect 16132 26812 18184 26840
rect 16132 26781 16160 26812
rect 14415 26744 14872 26772
rect 16117 26775 16175 26781
rect 14415 26741 14427 26744
rect 14369 26735 14427 26741
rect 16117 26741 16129 26775
rect 16163 26741 16175 26775
rect 16117 26735 16175 26741
rect 16758 26732 16764 26784
rect 16816 26772 16822 26784
rect 17497 26775 17555 26781
rect 17497 26772 17509 26775
rect 16816 26744 17509 26772
rect 16816 26732 16822 26744
rect 17497 26741 17509 26744
rect 17543 26741 17555 26775
rect 18156 26772 18184 26812
rect 19334 26800 19340 26852
rect 19392 26840 19398 26852
rect 21376 26840 21404 27016
rect 22370 27004 22376 27016
rect 22428 27004 22434 27056
rect 22002 26936 22008 26988
rect 22060 26936 22066 26988
rect 23400 26976 23428 27084
rect 23658 27072 23664 27124
rect 23716 27112 23722 27124
rect 25225 27115 25283 27121
rect 25225 27112 25237 27115
rect 23716 27084 25237 27112
rect 23716 27072 23722 27084
rect 25225 27081 25237 27084
rect 25271 27081 25283 27115
rect 25225 27075 25283 27081
rect 24305 27047 24363 27053
rect 24305 27013 24317 27047
rect 24351 27044 24363 27047
rect 24394 27044 24400 27056
rect 24351 27016 24400 27044
rect 24351 27013 24363 27016
rect 24305 27007 24363 27013
rect 24394 27004 24400 27016
rect 24452 27004 24458 27056
rect 23658 26976 23664 26988
rect 23400 26962 23664 26976
rect 23414 26948 23664 26962
rect 23658 26936 23664 26948
rect 23716 26936 23722 26988
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26976 24639 26979
rect 25222 26976 25228 26988
rect 24627 26948 25228 26976
rect 24627 26945 24639 26948
rect 24581 26939 24639 26945
rect 25222 26936 25228 26948
rect 25280 26936 25286 26988
rect 22281 26911 22339 26917
rect 22281 26877 22293 26911
rect 22327 26908 22339 26911
rect 25958 26908 25964 26920
rect 22327 26880 25964 26908
rect 22327 26877 22339 26880
rect 22281 26871 22339 26877
rect 25958 26868 25964 26880
rect 26016 26868 26022 26920
rect 19392 26812 21404 26840
rect 19392 26800 19398 26812
rect 18966 26772 18972 26784
rect 18156 26744 18972 26772
rect 17497 26735 17555 26741
rect 18966 26732 18972 26744
rect 19024 26732 19030 26784
rect 19058 26732 19064 26784
rect 19116 26772 19122 26784
rect 19797 26775 19855 26781
rect 19797 26772 19809 26775
rect 19116 26744 19809 26772
rect 19116 26732 19122 26744
rect 19797 26741 19809 26744
rect 19843 26741 19855 26775
rect 19797 26735 19855 26741
rect 20162 26732 20168 26784
rect 20220 26772 20226 26784
rect 20806 26772 20812 26784
rect 20220 26744 20812 26772
rect 20220 26732 20226 26744
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 21634 26732 21640 26784
rect 21692 26772 21698 26784
rect 23753 26775 23811 26781
rect 23753 26772 23765 26775
rect 21692 26744 23765 26772
rect 21692 26732 21698 26744
rect 23753 26741 23765 26744
rect 23799 26741 23811 26775
rect 23753 26735 23811 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8938 26568 8944 26580
rect 8619 26540 8944 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 8938 26528 8944 26540
rect 8996 26528 9002 26580
rect 9398 26528 9404 26580
rect 9456 26568 9462 26580
rect 10505 26571 10563 26577
rect 10505 26568 10517 26571
rect 9456 26540 10517 26568
rect 9456 26528 9462 26540
rect 10505 26537 10517 26540
rect 10551 26537 10563 26571
rect 13814 26568 13820 26580
rect 10505 26531 10563 26537
rect 10796 26540 13820 26568
rect 9125 26503 9183 26509
rect 9125 26469 9137 26503
rect 9171 26500 9183 26503
rect 10318 26500 10324 26512
rect 9171 26472 10324 26500
rect 9171 26469 9183 26472
rect 9125 26463 9183 26469
rect 6822 26324 6828 26376
rect 6880 26324 6886 26376
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 8478 26364 8484 26376
rect 7975 26336 8484 26364
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 8478 26324 8484 26336
rect 8536 26324 8542 26376
rect 9232 26373 9260 26472
rect 10318 26460 10324 26472
rect 10376 26460 10382 26512
rect 10594 26432 10600 26444
rect 9416 26404 10600 26432
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9217 26327 9275 26333
rect 7469 26299 7527 26305
rect 7469 26265 7481 26299
rect 7515 26296 7527 26299
rect 9416 26296 9444 26404
rect 10594 26392 10600 26404
rect 10652 26392 10658 26444
rect 9861 26367 9919 26373
rect 9861 26333 9873 26367
rect 9907 26364 9919 26367
rect 10796 26364 10824 26540
rect 13814 26528 13820 26540
rect 13872 26568 13878 26580
rect 14918 26568 14924 26580
rect 13872 26540 14924 26568
rect 13872 26528 13878 26540
rect 14918 26528 14924 26540
rect 14976 26528 14982 26580
rect 15102 26528 15108 26580
rect 15160 26568 15166 26580
rect 16301 26571 16359 26577
rect 16301 26568 16313 26571
rect 15160 26540 16313 26568
rect 15160 26528 15166 26540
rect 16301 26537 16313 26540
rect 16347 26537 16359 26571
rect 19334 26568 19340 26580
rect 16301 26531 16359 26537
rect 16592 26540 19340 26568
rect 12069 26503 12127 26509
rect 12069 26469 12081 26503
rect 12115 26500 12127 26503
rect 13446 26500 13452 26512
rect 12115 26472 13452 26500
rect 12115 26469 12127 26472
rect 12069 26463 12127 26469
rect 13446 26460 13452 26472
rect 13504 26460 13510 26512
rect 13541 26503 13599 26509
rect 13541 26469 13553 26503
rect 13587 26500 13599 26503
rect 13630 26500 13636 26512
rect 13587 26472 13636 26500
rect 13587 26469 13599 26472
rect 13541 26463 13599 26469
rect 13630 26460 13636 26472
rect 13688 26460 13694 26512
rect 14093 26503 14151 26509
rect 14093 26469 14105 26503
rect 14139 26500 14151 26503
rect 16592 26500 16620 26540
rect 19334 26528 19340 26540
rect 19392 26528 19398 26580
rect 19692 26571 19750 26577
rect 19692 26537 19704 26571
rect 19738 26568 19750 26571
rect 25130 26568 25136 26580
rect 19738 26540 25136 26568
rect 19738 26537 19750 26540
rect 19692 26531 19750 26537
rect 25130 26528 25136 26540
rect 25188 26528 25194 26580
rect 18322 26500 18328 26512
rect 14139 26472 16620 26500
rect 16684 26472 18328 26500
rect 14139 26469 14151 26472
rect 14093 26463 14151 26469
rect 11606 26392 11612 26444
rect 11664 26432 11670 26444
rect 12621 26435 12679 26441
rect 12621 26432 12633 26435
rect 11664 26404 12633 26432
rect 11664 26392 11670 26404
rect 12621 26401 12633 26404
rect 12667 26401 12679 26435
rect 12621 26395 12679 26401
rect 9907 26336 10824 26364
rect 9907 26333 9919 26336
rect 9861 26327 9919 26333
rect 10870 26324 10876 26376
rect 10928 26364 10934 26376
rect 10965 26367 11023 26373
rect 10965 26364 10977 26367
rect 10928 26336 10977 26364
rect 10928 26324 10934 26336
rect 10965 26333 10977 26336
rect 11011 26333 11023 26367
rect 12437 26367 12495 26373
rect 12437 26364 12449 26367
rect 10965 26327 11023 26333
rect 11072 26336 12449 26364
rect 7515 26268 9444 26296
rect 7515 26265 7527 26268
rect 7469 26259 7527 26265
rect 9490 26256 9496 26308
rect 9548 26296 9554 26308
rect 11072 26296 11100 26336
rect 12437 26333 12449 26336
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26364 12587 26367
rect 13538 26364 13544 26376
rect 12575 26336 13544 26364
rect 12575 26333 12587 26336
rect 12529 26327 12587 26333
rect 13538 26324 13544 26336
rect 13596 26324 13602 26376
rect 13725 26367 13783 26373
rect 13725 26333 13737 26367
rect 13771 26364 13783 26367
rect 14108 26364 14136 26463
rect 15010 26392 15016 26444
rect 15068 26392 15074 26444
rect 13771 26336 14136 26364
rect 15657 26367 15715 26373
rect 13771 26333 13783 26336
rect 13725 26327 13783 26333
rect 15657 26333 15669 26367
rect 15703 26364 15715 26367
rect 16684 26364 16712 26472
rect 18322 26460 18328 26472
rect 18380 26460 18386 26512
rect 21174 26460 21180 26512
rect 21232 26460 21238 26512
rect 24581 26503 24639 26509
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 25038 26500 25044 26512
rect 24627 26472 25044 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 25038 26460 25044 26472
rect 25096 26460 25102 26512
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 19429 26435 19487 26441
rect 19429 26432 19441 26435
rect 17920 26404 19441 26432
rect 17920 26392 17926 26404
rect 19429 26401 19441 26404
rect 19475 26432 19487 26435
rect 19702 26432 19708 26444
rect 19475 26404 19708 26432
rect 19475 26401 19487 26404
rect 19429 26395 19487 26401
rect 19702 26392 19708 26404
rect 19760 26432 19766 26444
rect 20438 26432 20444 26444
rect 19760 26404 20444 26432
rect 19760 26392 19766 26404
rect 20438 26392 20444 26404
rect 20496 26392 20502 26444
rect 21358 26392 21364 26444
rect 21416 26432 21422 26444
rect 21910 26432 21916 26444
rect 21416 26404 21916 26432
rect 21416 26392 21422 26404
rect 21910 26392 21916 26404
rect 21968 26392 21974 26444
rect 22002 26392 22008 26444
rect 22060 26432 22066 26444
rect 22281 26435 22339 26441
rect 22281 26432 22293 26435
rect 22060 26404 22293 26432
rect 22060 26392 22066 26404
rect 22281 26401 22293 26404
rect 22327 26432 22339 26435
rect 23290 26432 23296 26444
rect 22327 26404 23296 26432
rect 22327 26401 22339 26404
rect 22281 26395 22339 26401
rect 23290 26392 23296 26404
rect 23348 26392 23354 26444
rect 24029 26435 24087 26441
rect 24029 26401 24041 26435
rect 24075 26432 24087 26435
rect 24302 26432 24308 26444
rect 24075 26404 24308 26432
rect 24075 26401 24087 26404
rect 24029 26395 24087 26401
rect 24302 26392 24308 26404
rect 24360 26392 24366 26444
rect 25225 26435 25283 26441
rect 25225 26401 25237 26435
rect 25271 26432 25283 26435
rect 25314 26432 25320 26444
rect 25271 26404 25320 26432
rect 25271 26401 25283 26404
rect 25225 26395 25283 26401
rect 25314 26392 25320 26404
rect 25372 26392 25378 26444
rect 15703 26336 16712 26364
rect 15703 26333 15715 26336
rect 15657 26327 15715 26333
rect 16758 26324 16764 26376
rect 16816 26324 16822 26376
rect 17957 26367 18015 26373
rect 17957 26333 17969 26367
rect 18003 26364 18015 26367
rect 18690 26364 18696 26376
rect 18003 26336 18696 26364
rect 18003 26333 18015 26336
rect 17957 26327 18015 26333
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 18782 26324 18788 26376
rect 18840 26364 18846 26376
rect 18966 26364 18972 26376
rect 18840 26336 18972 26364
rect 18840 26324 18846 26336
rect 18966 26324 18972 26336
rect 19024 26324 19030 26376
rect 20806 26324 20812 26376
rect 20864 26364 20870 26376
rect 20864 26336 21956 26364
rect 20864 26324 20870 26336
rect 9548 26268 11100 26296
rect 9548 26256 9554 26268
rect 11514 26256 11520 26308
rect 11572 26296 11578 26308
rect 11609 26299 11667 26305
rect 11609 26296 11621 26299
rect 11572 26268 11621 26296
rect 11572 26256 11578 26268
rect 11609 26265 11621 26268
rect 11655 26265 11667 26299
rect 14829 26299 14887 26305
rect 11609 26259 11667 26265
rect 12406 26268 14504 26296
rect 12406 26240 12434 26268
rect 12342 26188 12348 26240
rect 12400 26200 12434 26240
rect 12400 26188 12406 26200
rect 13538 26188 13544 26240
rect 13596 26228 13602 26240
rect 13722 26228 13728 26240
rect 13596 26200 13728 26228
rect 13596 26188 13602 26200
rect 13722 26188 13728 26200
rect 13780 26188 13786 26240
rect 14476 26237 14504 26268
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 14875 26268 15148 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 14461 26231 14519 26237
rect 14461 26197 14473 26231
rect 14507 26197 14519 26231
rect 14461 26191 14519 26197
rect 14918 26188 14924 26240
rect 14976 26188 14982 26240
rect 15120 26228 15148 26268
rect 15194 26256 15200 26308
rect 15252 26296 15258 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 15252 26268 17417 26296
rect 15252 26256 15258 26268
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17405 26259 17463 26265
rect 18414 26256 18420 26308
rect 18472 26296 18478 26308
rect 21637 26299 21695 26305
rect 21637 26296 21649 26299
rect 18472 26268 20116 26296
rect 18472 26256 18478 26268
rect 15746 26228 15752 26240
rect 15120 26200 15752 26228
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 18598 26188 18604 26240
rect 18656 26188 18662 26240
rect 20088 26228 20116 26268
rect 21008 26268 21649 26296
rect 21008 26228 21036 26268
rect 21637 26265 21649 26268
rect 21683 26265 21695 26299
rect 21637 26259 21695 26265
rect 20088 26200 21036 26228
rect 21928 26228 21956 26336
rect 23658 26324 23664 26376
rect 23716 26324 23722 26376
rect 24394 26324 24400 26376
rect 24452 26364 24458 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 24452 26336 24961 26364
rect 24452 26324 24458 26336
rect 24949 26333 24961 26336
rect 24995 26333 25007 26367
rect 24949 26327 25007 26333
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26364 25099 26367
rect 25406 26364 25412 26376
rect 25087 26336 25412 26364
rect 25087 26333 25099 26336
rect 25041 26327 25099 26333
rect 22002 26256 22008 26308
rect 22060 26296 22066 26308
rect 22557 26299 22615 26305
rect 22557 26296 22569 26299
rect 22060 26268 22569 26296
rect 22060 26256 22066 26268
rect 22557 26265 22569 26268
rect 22603 26265 22615 26299
rect 24964 26296 24992 26327
rect 25406 26324 25412 26336
rect 25464 26324 25470 26376
rect 25774 26296 25780 26308
rect 24964 26268 25780 26296
rect 22557 26259 22615 26265
rect 25774 26256 25780 26268
rect 25832 26256 25838 26308
rect 22094 26228 22100 26240
rect 21928 26200 22100 26228
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 9508 25996 11008 26024
rect 9508 25956 9536 25996
rect 10980 25968 11008 25996
rect 11330 25984 11336 26036
rect 11388 26024 11394 26036
rect 12618 26024 12624 26036
rect 11388 25996 12624 26024
rect 11388 25984 11394 25996
rect 12618 25984 12624 25996
rect 12676 26024 12682 26036
rect 12676 25996 12940 26024
rect 12676 25984 12682 25996
rect 9416 25928 9536 25956
rect 9416 25897 9444 25928
rect 9674 25916 9680 25968
rect 9732 25916 9738 25968
rect 10962 25916 10968 25968
rect 11020 25956 11026 25968
rect 12526 25956 12532 25968
rect 11020 25928 12532 25956
rect 11020 25916 11026 25928
rect 12526 25916 12532 25928
rect 12584 25956 12590 25968
rect 12912 25956 12940 25996
rect 13722 25984 13728 26036
rect 13780 26024 13786 26036
rect 13780 25996 14412 26024
rect 13780 25984 13786 25996
rect 14384 25956 14412 25996
rect 15378 25984 15384 26036
rect 15436 25984 15442 26036
rect 15473 26027 15531 26033
rect 15473 25993 15485 26027
rect 15519 26024 15531 26027
rect 16666 26024 16672 26036
rect 15519 25996 16672 26024
rect 15519 25993 15531 25996
rect 15473 25987 15531 25993
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 17221 26027 17279 26033
rect 17221 25993 17233 26027
rect 17267 26024 17279 26027
rect 17586 26024 17592 26036
rect 17267 25996 17592 26024
rect 17267 25993 17279 25996
rect 17221 25987 17279 25993
rect 17586 25984 17592 25996
rect 17644 25984 17650 26036
rect 18414 25984 18420 26036
rect 18472 25984 18478 26036
rect 18509 26027 18567 26033
rect 18509 25993 18521 26027
rect 18555 26024 18567 26027
rect 20622 26024 20628 26036
rect 18555 25996 20628 26024
rect 18555 25993 18567 25996
rect 18509 25987 18567 25993
rect 20622 25984 20628 25996
rect 20680 25984 20686 26036
rect 21266 25984 21272 26036
rect 21324 25984 21330 26036
rect 21542 25984 21548 26036
rect 21600 25984 21606 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 24118 26024 24124 26036
rect 22152 25996 24124 26024
rect 22152 25984 22158 25996
rect 24118 25984 24124 25996
rect 24176 25984 24182 26036
rect 17604 25956 17632 25984
rect 19061 25959 19119 25965
rect 19061 25956 19073 25959
rect 12584 25928 12848 25956
rect 12912 25928 13570 25956
rect 14384 25928 17448 25956
rect 17604 25928 19073 25956
rect 12584 25916 12590 25928
rect 7193 25891 7251 25897
rect 7193 25857 7205 25891
rect 7239 25857 7251 25891
rect 7193 25851 7251 25857
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25857 8355 25891
rect 8297 25851 8355 25857
rect 9401 25891 9459 25897
rect 9401 25857 9413 25891
rect 9447 25857 9459 25891
rect 9401 25851 9459 25857
rect 7208 25752 7236 25851
rect 8312 25820 8340 25851
rect 10778 25848 10784 25900
rect 10836 25888 10842 25900
rect 11330 25888 11336 25900
rect 10836 25860 11336 25888
rect 10836 25848 10842 25860
rect 11330 25848 11336 25860
rect 11388 25848 11394 25900
rect 11606 25848 11612 25900
rect 11664 25888 11670 25900
rect 12820 25897 12848 25928
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 11664 25860 11713 25888
rect 11664 25848 11670 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 12805 25891 12863 25897
rect 12805 25857 12817 25891
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 14918 25848 14924 25900
rect 14976 25888 14982 25900
rect 15102 25888 15108 25900
rect 14976 25860 15108 25888
rect 14976 25848 14982 25860
rect 15102 25848 15108 25860
rect 15160 25888 15166 25900
rect 15160 25860 15700 25888
rect 15160 25848 15166 25860
rect 10318 25820 10324 25832
rect 8312 25792 10324 25820
rect 10318 25780 10324 25792
rect 10376 25780 10382 25832
rect 10686 25780 10692 25832
rect 10744 25820 10750 25832
rect 12345 25823 12403 25829
rect 12345 25820 12357 25823
rect 10744 25792 12357 25820
rect 10744 25780 10750 25792
rect 12345 25789 12357 25792
rect 12391 25789 12403 25823
rect 12345 25783 12403 25789
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25820 13139 25823
rect 15470 25820 15476 25832
rect 13127 25792 15476 25820
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 15470 25780 15476 25792
rect 15528 25780 15534 25832
rect 15565 25823 15623 25829
rect 15565 25789 15577 25823
rect 15611 25789 15623 25823
rect 15672 25820 15700 25860
rect 16114 25848 16120 25900
rect 16172 25888 16178 25900
rect 16172 25860 17356 25888
rect 16172 25848 16178 25860
rect 16301 25823 16359 25829
rect 16301 25820 16313 25823
rect 15672 25792 16313 25820
rect 15565 25783 15623 25789
rect 16301 25789 16313 25792
rect 16347 25820 16359 25823
rect 16666 25820 16672 25832
rect 16347 25792 16672 25820
rect 16347 25789 16359 25792
rect 16301 25783 16359 25789
rect 12802 25752 12808 25764
rect 7208 25724 9076 25752
rect 9048 25696 9076 25724
rect 11164 25724 12808 25752
rect 7466 25644 7472 25696
rect 7524 25684 7530 25696
rect 7837 25687 7895 25693
rect 7837 25684 7849 25687
rect 7524 25656 7849 25684
rect 7524 25644 7530 25656
rect 7837 25653 7849 25656
rect 7883 25653 7895 25687
rect 7837 25647 7895 25653
rect 8938 25644 8944 25696
rect 8996 25644 9002 25696
rect 9030 25644 9036 25696
rect 9088 25684 9094 25696
rect 11164 25693 11192 25724
rect 12802 25712 12808 25724
rect 12860 25712 12866 25764
rect 15580 25752 15608 25783
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 17328 25829 17356 25860
rect 17420 25829 17448 25928
rect 19061 25925 19073 25928
rect 19107 25925 19119 25959
rect 21560 25956 21588 25984
rect 23290 25956 23296 25968
rect 19061 25919 19119 25925
rect 19168 25928 21588 25956
rect 23124 25928 23296 25956
rect 18782 25888 18788 25900
rect 17512 25860 18788 25888
rect 17313 25823 17371 25829
rect 17313 25789 17325 25823
rect 17359 25789 17371 25823
rect 17313 25783 17371 25789
rect 17405 25823 17463 25829
rect 17405 25789 17417 25823
rect 17451 25789 17463 25823
rect 17405 25783 17463 25789
rect 14568 25724 15608 25752
rect 11149 25687 11207 25693
rect 11149 25684 11161 25687
rect 9088 25656 11161 25684
rect 9088 25644 9094 25656
rect 11149 25653 11161 25656
rect 11195 25653 11207 25687
rect 11149 25647 11207 25653
rect 11698 25644 11704 25696
rect 11756 25684 11762 25696
rect 14568 25693 14596 25724
rect 15746 25712 15752 25764
rect 15804 25752 15810 25764
rect 16393 25755 16451 25761
rect 16393 25752 16405 25755
rect 15804 25724 16405 25752
rect 15804 25712 15810 25724
rect 16393 25721 16405 25724
rect 16439 25721 16451 25755
rect 17328 25752 17356 25783
rect 17512 25752 17540 25860
rect 18782 25848 18788 25860
rect 18840 25888 18846 25900
rect 19168 25888 19196 25928
rect 18840 25860 19196 25888
rect 18840 25848 18846 25860
rect 19518 25848 19524 25900
rect 19576 25848 19582 25900
rect 20165 25891 20223 25897
rect 20165 25857 20177 25891
rect 20211 25888 20223 25891
rect 20625 25891 20683 25897
rect 20625 25888 20637 25891
rect 20211 25860 20637 25888
rect 20211 25857 20223 25860
rect 20165 25851 20223 25857
rect 20625 25857 20637 25860
rect 20671 25857 20683 25891
rect 20625 25851 20683 25857
rect 21542 25848 21548 25900
rect 21600 25888 21606 25900
rect 23124 25897 23152 25928
rect 23290 25916 23296 25928
rect 23348 25916 23354 25968
rect 23382 25916 23388 25968
rect 23440 25916 23446 25968
rect 23658 25916 23664 25968
rect 23716 25956 23722 25968
rect 23716 25928 23874 25956
rect 23716 25916 23722 25928
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21600 25860 22017 25888
rect 21600 25848 21606 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 23109 25891 23167 25897
rect 23109 25857 23121 25891
rect 23155 25857 23167 25891
rect 23109 25851 23167 25857
rect 18693 25823 18751 25829
rect 18693 25789 18705 25823
rect 18739 25820 18751 25823
rect 18874 25820 18880 25832
rect 18739 25792 18880 25820
rect 18739 25789 18751 25792
rect 18693 25783 18751 25789
rect 18874 25780 18880 25792
rect 18932 25780 18938 25832
rect 23382 25780 23388 25832
rect 23440 25820 23446 25832
rect 24857 25823 24915 25829
rect 24857 25820 24869 25823
rect 23440 25792 24869 25820
rect 23440 25780 23446 25792
rect 24857 25789 24869 25792
rect 24903 25789 24915 25823
rect 24857 25783 24915 25789
rect 17328 25724 17540 25752
rect 16393 25715 16451 25721
rect 18046 25712 18052 25764
rect 18104 25712 18110 25764
rect 14553 25687 14611 25693
rect 14553 25684 14565 25687
rect 11756 25656 14565 25684
rect 11756 25644 11762 25656
rect 14553 25653 14565 25656
rect 14599 25653 14611 25687
rect 14553 25647 14611 25653
rect 14734 25644 14740 25696
rect 14792 25684 14798 25696
rect 15013 25687 15071 25693
rect 15013 25684 15025 25687
rect 14792 25656 15025 25684
rect 14792 25644 14798 25656
rect 15013 25653 15025 25656
rect 15059 25653 15071 25687
rect 15013 25647 15071 25653
rect 15378 25644 15384 25696
rect 15436 25684 15442 25696
rect 16482 25684 16488 25696
rect 15436 25656 16488 25684
rect 15436 25644 15442 25656
rect 16482 25644 16488 25656
rect 16540 25644 16546 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 16853 25687 16911 25693
rect 16853 25684 16865 25687
rect 16632 25656 16865 25684
rect 16632 25644 16638 25656
rect 16853 25653 16865 25656
rect 16899 25653 16911 25687
rect 16853 25647 16911 25653
rect 22649 25687 22707 25693
rect 22649 25653 22661 25687
rect 22695 25684 22707 25687
rect 24578 25684 24584 25696
rect 22695 25656 24584 25684
rect 22695 25653 22707 25656
rect 22649 25647 22707 25653
rect 24578 25644 24584 25656
rect 24636 25644 24642 25696
rect 25222 25644 25228 25696
rect 25280 25644 25286 25696
rect 25406 25644 25412 25696
rect 25464 25644 25470 25696
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 9382 25483 9440 25489
rect 9382 25480 9394 25483
rect 8996 25452 9394 25480
rect 8996 25440 9002 25452
rect 9382 25449 9394 25452
rect 9428 25449 9440 25483
rect 9382 25443 9440 25449
rect 10134 25440 10140 25492
rect 10192 25480 10198 25492
rect 10594 25480 10600 25492
rect 10192 25452 10600 25480
rect 10192 25440 10198 25452
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 10873 25483 10931 25489
rect 10873 25449 10885 25483
rect 10919 25480 10931 25483
rect 10919 25452 12664 25480
rect 10919 25449 10931 25452
rect 10873 25443 10931 25449
rect 10502 25372 10508 25424
rect 10560 25412 10566 25424
rect 10888 25412 10916 25443
rect 10560 25384 10916 25412
rect 12636 25412 12664 25452
rect 13538 25440 13544 25492
rect 13596 25440 13602 25492
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 14507 25452 17540 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 12636 25384 14596 25412
rect 10560 25372 10566 25384
rect 9125 25347 9183 25353
rect 9125 25313 9137 25347
rect 9171 25344 9183 25347
rect 10962 25344 10968 25356
rect 9171 25316 10968 25344
rect 9171 25313 9183 25316
rect 9125 25307 9183 25313
rect 10962 25304 10968 25316
rect 11020 25344 11026 25356
rect 11333 25347 11391 25353
rect 11333 25344 11345 25347
rect 11020 25316 11345 25344
rect 11020 25304 11026 25316
rect 11333 25313 11345 25316
rect 11379 25313 11391 25347
rect 11333 25307 11391 25313
rect 11609 25347 11667 25353
rect 11609 25313 11621 25347
rect 11655 25344 11667 25347
rect 14458 25344 14464 25356
rect 11655 25316 14464 25344
rect 11655 25313 11667 25316
rect 11609 25307 11667 25313
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 7929 25279 7987 25285
rect 7929 25245 7941 25279
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 7944 25208 7972 25239
rect 13446 25236 13452 25288
rect 13504 25276 13510 25288
rect 13725 25279 13783 25285
rect 13725 25276 13737 25279
rect 13504 25248 13737 25276
rect 13504 25236 13510 25248
rect 13725 25245 13737 25248
rect 13771 25245 13783 25279
rect 14568 25276 14596 25384
rect 14642 25372 14648 25424
rect 14700 25412 14706 25424
rect 14700 25384 15056 25412
rect 14700 25372 14706 25384
rect 14826 25304 14832 25356
rect 14884 25344 14890 25356
rect 15028 25353 15056 25384
rect 14921 25347 14979 25353
rect 14921 25344 14933 25347
rect 14884 25316 14933 25344
rect 14884 25304 14890 25316
rect 14921 25313 14933 25316
rect 14967 25313 14979 25347
rect 14921 25307 14979 25313
rect 15013 25347 15071 25353
rect 15013 25313 15025 25347
rect 15059 25313 15071 25347
rect 15013 25307 15071 25313
rect 15562 25304 15568 25356
rect 15620 25344 15626 25356
rect 16209 25347 16267 25353
rect 16209 25344 16221 25347
rect 15620 25316 16221 25344
rect 15620 25304 15626 25316
rect 16209 25313 16221 25316
rect 16255 25313 16267 25347
rect 17512 25344 17540 25452
rect 18690 25440 18696 25492
rect 18748 25440 18754 25492
rect 19061 25483 19119 25489
rect 19061 25449 19073 25483
rect 19107 25480 19119 25483
rect 19150 25480 19156 25492
rect 19107 25452 19156 25480
rect 19107 25449 19119 25452
rect 19061 25443 19119 25449
rect 19150 25440 19156 25452
rect 19208 25440 19214 25492
rect 19518 25440 19524 25492
rect 19576 25480 19582 25492
rect 20165 25483 20223 25489
rect 20165 25480 20177 25483
rect 19576 25452 20177 25480
rect 19576 25440 19582 25452
rect 20165 25449 20177 25452
rect 20211 25449 20223 25483
rect 20165 25443 20223 25449
rect 20714 25440 20720 25492
rect 20772 25480 20778 25492
rect 21910 25480 21916 25492
rect 20772 25452 21916 25480
rect 20772 25440 20778 25452
rect 21910 25440 21916 25452
rect 21968 25440 21974 25492
rect 25225 25483 25283 25489
rect 25225 25449 25237 25483
rect 25271 25480 25283 25483
rect 25682 25480 25688 25492
rect 25271 25452 25688 25480
rect 25271 25449 25283 25452
rect 25225 25443 25283 25449
rect 25682 25440 25688 25452
rect 25740 25440 25746 25492
rect 17589 25415 17647 25421
rect 17589 25381 17601 25415
rect 17635 25412 17647 25415
rect 24118 25412 24124 25424
rect 17635 25384 24124 25412
rect 17635 25381 17647 25384
rect 17589 25375 17647 25381
rect 24118 25372 24124 25384
rect 24176 25372 24182 25424
rect 17512 25316 20944 25344
rect 16209 25307 16267 25313
rect 14568 25248 15056 25276
rect 13725 25239 13783 25245
rect 15028 25220 15056 25248
rect 16114 25236 16120 25288
rect 16172 25236 16178 25288
rect 16945 25279 17003 25285
rect 16945 25245 16957 25279
rect 16991 25276 17003 25279
rect 17586 25276 17592 25288
rect 16991 25248 17592 25276
rect 16991 25245 17003 25248
rect 16945 25239 17003 25245
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 18049 25279 18107 25285
rect 18049 25245 18061 25279
rect 18095 25276 18107 25279
rect 19058 25276 19064 25288
rect 18095 25248 19064 25276
rect 18095 25245 18107 25248
rect 18049 25239 18107 25245
rect 19058 25236 19064 25248
rect 19116 25236 19122 25288
rect 19521 25279 19579 25285
rect 19521 25245 19533 25279
rect 19567 25245 19579 25279
rect 19521 25239 19579 25245
rect 9674 25208 9680 25220
rect 7944 25180 9680 25208
rect 9674 25168 9680 25180
rect 9732 25168 9738 25220
rect 10778 25208 10784 25220
rect 10626 25180 10784 25208
rect 10778 25168 10784 25180
rect 10836 25168 10842 25220
rect 12618 25168 12624 25220
rect 12676 25168 12682 25220
rect 13814 25208 13820 25220
rect 13096 25180 13820 25208
rect 8573 25143 8631 25149
rect 8573 25109 8585 25143
rect 8619 25140 8631 25143
rect 10134 25140 10140 25152
rect 8619 25112 10140 25140
rect 8619 25109 8631 25112
rect 8573 25103 8631 25109
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 13096 25149 13124 25180
rect 13814 25168 13820 25180
rect 13872 25168 13878 25220
rect 14182 25168 14188 25220
rect 14240 25208 14246 25220
rect 14829 25211 14887 25217
rect 14829 25208 14841 25211
rect 14240 25180 14841 25208
rect 14240 25168 14246 25180
rect 14829 25177 14841 25180
rect 14875 25177 14887 25211
rect 14829 25171 14887 25177
rect 15010 25168 15016 25220
rect 15068 25168 15074 25220
rect 16758 25168 16764 25220
rect 16816 25208 16822 25220
rect 18506 25208 18512 25220
rect 16816 25180 18512 25208
rect 16816 25168 16822 25180
rect 18506 25168 18512 25180
rect 18564 25168 18570 25220
rect 19536 25208 19564 25239
rect 20714 25236 20720 25288
rect 20772 25236 20778 25288
rect 20916 25276 20944 25316
rect 20990 25304 20996 25356
rect 21048 25344 21054 25356
rect 22005 25347 22063 25353
rect 22005 25344 22017 25347
rect 21048 25316 22017 25344
rect 21048 25304 21054 25316
rect 22005 25313 22017 25316
rect 22051 25313 22063 25347
rect 22005 25307 22063 25313
rect 21450 25276 21456 25288
rect 20916 25248 21456 25276
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 21910 25236 21916 25288
rect 21968 25236 21974 25288
rect 22554 25236 22560 25288
rect 22612 25276 22618 25288
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 22612 25248 22661 25276
rect 22612 25236 22618 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 24394 25236 24400 25288
rect 24452 25276 24458 25288
rect 24581 25279 24639 25285
rect 24581 25276 24593 25279
rect 24452 25248 24593 25276
rect 24452 25236 24458 25248
rect 24581 25245 24593 25248
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 21174 25208 21180 25220
rect 19536 25180 21180 25208
rect 21174 25168 21180 25180
rect 21232 25168 21238 25220
rect 22830 25168 22836 25220
rect 22888 25168 22894 25220
rect 23845 25211 23903 25217
rect 23845 25177 23857 25211
rect 23891 25208 23903 25211
rect 24946 25208 24952 25220
rect 23891 25180 24952 25208
rect 23891 25177 23903 25180
rect 23845 25171 23903 25177
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 13081 25143 13139 25149
rect 13081 25109 13093 25143
rect 13127 25109 13139 25143
rect 13081 25103 13139 25109
rect 13170 25100 13176 25152
rect 13228 25140 13234 25152
rect 13906 25140 13912 25152
rect 13228 25112 13912 25140
rect 13228 25100 13234 25112
rect 13906 25100 13912 25112
rect 13964 25100 13970 25152
rect 14642 25100 14648 25152
rect 14700 25140 14706 25152
rect 15657 25143 15715 25149
rect 15657 25140 15669 25143
rect 14700 25112 15669 25140
rect 14700 25100 14706 25112
rect 15657 25109 15669 25112
rect 15703 25109 15715 25143
rect 15657 25103 15715 25109
rect 16022 25100 16028 25152
rect 16080 25100 16086 25152
rect 16390 25100 16396 25152
rect 16448 25140 16454 25152
rect 18322 25140 18328 25152
rect 16448 25112 18328 25140
rect 16448 25100 16454 25112
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 20806 25100 20812 25152
rect 20864 25100 20870 25152
rect 20898 25100 20904 25152
rect 20956 25140 20962 25152
rect 21453 25143 21511 25149
rect 21453 25140 21465 25143
rect 20956 25112 21465 25140
rect 20956 25100 20962 25112
rect 21453 25109 21465 25112
rect 21499 25109 21511 25143
rect 21453 25103 21511 25109
rect 21821 25143 21879 25149
rect 21821 25109 21833 25143
rect 21867 25140 21879 25143
rect 21910 25140 21916 25152
rect 21867 25112 21916 25140
rect 21867 25109 21879 25112
rect 21821 25103 21879 25109
rect 21910 25100 21916 25112
rect 21968 25100 21974 25152
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 22848 25140 22876 25168
rect 22612 25112 22876 25140
rect 22612 25100 22618 25112
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 9582 24896 9588 24948
rect 9640 24936 9646 24948
rect 10502 24936 10508 24948
rect 9640 24908 10508 24936
rect 9640 24896 9646 24908
rect 10502 24896 10508 24908
rect 10560 24896 10566 24948
rect 14461 24939 14519 24945
rect 14461 24905 14473 24939
rect 14507 24936 14519 24939
rect 15378 24936 15384 24948
rect 14507 24908 15384 24936
rect 14507 24905 14519 24908
rect 14461 24899 14519 24905
rect 15378 24896 15384 24908
rect 15436 24896 15442 24948
rect 16114 24896 16120 24948
rect 16172 24936 16178 24948
rect 16298 24936 16304 24948
rect 16172 24908 16304 24936
rect 16172 24896 16178 24908
rect 16298 24896 16304 24908
rect 16356 24936 16362 24948
rect 16393 24939 16451 24945
rect 16393 24936 16405 24939
rect 16356 24908 16405 24936
rect 16356 24896 16362 24908
rect 16393 24905 16405 24908
rect 16439 24905 16451 24939
rect 16393 24899 16451 24905
rect 16482 24896 16488 24948
rect 16540 24936 16546 24948
rect 17221 24939 17279 24945
rect 17221 24936 17233 24939
rect 16540 24908 17233 24936
rect 16540 24896 16546 24908
rect 17221 24905 17233 24908
rect 17267 24905 17279 24939
rect 17221 24899 17279 24905
rect 17313 24939 17371 24945
rect 17313 24905 17325 24939
rect 17359 24936 17371 24939
rect 17494 24936 17500 24948
rect 17359 24908 17500 24936
rect 17359 24905 17371 24908
rect 17313 24899 17371 24905
rect 17494 24896 17500 24908
rect 17552 24936 17558 24948
rect 17552 24908 17632 24936
rect 17552 24896 17558 24908
rect 10778 24868 10784 24880
rect 10074 24840 10784 24868
rect 10778 24828 10784 24840
rect 10836 24828 10842 24880
rect 12802 24828 12808 24880
rect 12860 24868 12866 24880
rect 12860 24840 13400 24868
rect 12860 24828 12866 24840
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 8570 24760 8576 24812
rect 8628 24760 8634 24812
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 13170 24760 13176 24812
rect 13228 24760 13234 24812
rect 13262 24760 13268 24812
rect 13320 24760 13326 24812
rect 13372 24741 13400 24840
rect 13538 24828 13544 24880
rect 13596 24868 13602 24880
rect 13722 24868 13728 24880
rect 13596 24840 13728 24868
rect 13596 24828 13602 24840
rect 13722 24828 13728 24840
rect 13780 24828 13786 24880
rect 14369 24871 14427 24877
rect 14369 24837 14381 24871
rect 14415 24868 14427 24871
rect 15654 24868 15660 24880
rect 14415 24840 15660 24868
rect 14415 24837 14427 24840
rect 14369 24831 14427 24837
rect 15654 24828 15660 24840
rect 15712 24828 15718 24880
rect 17604 24868 17632 24908
rect 17678 24896 17684 24948
rect 17736 24936 17742 24948
rect 17865 24939 17923 24945
rect 17865 24936 17877 24939
rect 17736 24908 17877 24936
rect 17736 24896 17742 24908
rect 17865 24905 17877 24908
rect 17911 24936 17923 24939
rect 18598 24936 18604 24948
rect 17911 24908 18604 24936
rect 17911 24905 17923 24908
rect 17865 24899 17923 24905
rect 18598 24896 18604 24908
rect 18656 24896 18662 24948
rect 19150 24936 19156 24948
rect 18708 24908 19156 24936
rect 18708 24880 18736 24908
rect 19150 24896 19156 24908
rect 19208 24896 19214 24948
rect 20714 24896 20720 24948
rect 20772 24936 20778 24948
rect 21821 24939 21879 24945
rect 21821 24936 21833 24939
rect 20772 24908 21833 24936
rect 20772 24896 20778 24908
rect 21821 24905 21833 24908
rect 21867 24905 21879 24939
rect 21821 24899 21879 24905
rect 22741 24939 22799 24945
rect 22741 24905 22753 24939
rect 22787 24936 22799 24939
rect 24026 24936 24032 24948
rect 22787 24908 24032 24936
rect 22787 24905 22799 24908
rect 22741 24899 22799 24905
rect 24026 24896 24032 24908
rect 24084 24896 24090 24948
rect 18690 24868 18696 24880
rect 17144 24840 17356 24868
rect 17604 24840 18696 24868
rect 15194 24760 15200 24812
rect 15252 24760 15258 24812
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 15841 24803 15899 24809
rect 15841 24800 15853 24803
rect 15528 24772 15853 24800
rect 15528 24760 15534 24772
rect 15841 24769 15853 24772
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 16206 24760 16212 24812
rect 16264 24800 16270 24812
rect 17144 24800 17172 24840
rect 16264 24772 17172 24800
rect 17328 24800 17356 24840
rect 18690 24828 18696 24840
rect 18748 24828 18754 24880
rect 18877 24871 18935 24877
rect 18877 24837 18889 24871
rect 18923 24868 18935 24871
rect 19978 24868 19984 24880
rect 18923 24840 19984 24868
rect 18923 24837 18935 24840
rect 18877 24831 18935 24837
rect 19978 24828 19984 24840
rect 20036 24828 20042 24880
rect 21910 24868 21916 24880
rect 21206 24840 21916 24868
rect 21910 24828 21916 24840
rect 21968 24828 21974 24880
rect 25222 24868 25228 24880
rect 25070 24840 25228 24868
rect 25222 24828 25228 24840
rect 25280 24828 25286 24880
rect 17328 24772 17448 24800
rect 16264 24760 16270 24772
rect 8113 24735 8171 24741
rect 8113 24701 8125 24735
rect 8159 24732 8171 24735
rect 8849 24735 8907 24741
rect 8849 24732 8861 24735
rect 8159 24704 8861 24732
rect 8159 24701 8171 24704
rect 8113 24695 8171 24701
rect 8849 24701 8861 24704
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 13357 24735 13415 24741
rect 13357 24701 13369 24735
rect 13403 24701 13415 24735
rect 13357 24695 13415 24701
rect 14645 24735 14703 24741
rect 14645 24701 14657 24735
rect 14691 24732 14703 24735
rect 15010 24732 15016 24744
rect 14691 24704 15016 24732
rect 14691 24701 14703 24704
rect 14645 24695 14703 24701
rect 10980 24664 11008 24695
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 16482 24692 16488 24744
rect 16540 24732 16546 24744
rect 17310 24732 17316 24744
rect 16540 24704 17316 24732
rect 16540 24692 16546 24704
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 17420 24741 17448 24772
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19702 24800 19708 24812
rect 19392 24772 19708 24800
rect 19392 24760 19398 24772
rect 19702 24760 19708 24772
rect 19760 24760 19766 24812
rect 21266 24760 21272 24812
rect 21324 24800 21330 24812
rect 21324 24772 22508 24800
rect 21324 24760 21330 24772
rect 17405 24735 17463 24741
rect 17405 24701 17417 24735
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 18141 24735 18199 24741
rect 18141 24701 18153 24735
rect 18187 24732 18199 24735
rect 18322 24732 18328 24744
rect 18187 24704 18328 24732
rect 18187 24701 18199 24704
rect 18141 24695 18199 24701
rect 18322 24692 18328 24704
rect 18380 24692 18386 24744
rect 18969 24735 19027 24741
rect 18969 24701 18981 24735
rect 19015 24701 19027 24735
rect 18969 24695 19027 24701
rect 18414 24664 18420 24676
rect 10980 24636 14504 24664
rect 9858 24556 9864 24608
rect 9916 24596 9922 24608
rect 10321 24599 10379 24605
rect 10321 24596 10333 24599
rect 9916 24568 10333 24596
rect 9916 24556 9922 24568
rect 10321 24565 10333 24568
rect 10367 24596 10379 24599
rect 10686 24596 10692 24608
rect 10367 24568 10692 24596
rect 10367 24565 10379 24568
rect 10321 24559 10379 24565
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 10870 24556 10876 24608
rect 10928 24596 10934 24608
rect 12345 24599 12403 24605
rect 12345 24596 12357 24599
rect 10928 24568 12357 24596
rect 10928 24556 10934 24568
rect 12345 24565 12357 24568
rect 12391 24565 12403 24599
rect 12345 24559 12403 24565
rect 12526 24556 12532 24608
rect 12584 24596 12590 24608
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12584 24568 12817 24596
rect 12584 24556 12590 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 12805 24559 12863 24565
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 14001 24599 14059 24605
rect 14001 24596 14013 24599
rect 13412 24568 14013 24596
rect 13412 24556 13418 24568
rect 14001 24565 14013 24568
rect 14047 24565 14059 24599
rect 14476 24596 14504 24636
rect 14660 24636 18420 24664
rect 14660 24596 14688 24636
rect 18414 24624 18420 24636
rect 18472 24624 18478 24676
rect 18506 24624 18512 24676
rect 18564 24624 18570 24676
rect 14476 24568 14688 24596
rect 16209 24599 16267 24605
rect 14001 24559 14059 24565
rect 16209 24565 16221 24599
rect 16255 24596 16267 24599
rect 16482 24596 16488 24608
rect 16255 24568 16488 24596
rect 16255 24565 16267 24568
rect 16209 24559 16267 24565
rect 16482 24556 16488 24568
rect 16540 24556 16546 24608
rect 16853 24599 16911 24605
rect 16853 24565 16865 24599
rect 16899 24596 16911 24599
rect 16942 24596 16948 24608
rect 16899 24568 16948 24596
rect 16899 24565 16911 24568
rect 16853 24559 16911 24565
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 18984 24596 19012 24695
rect 19058 24692 19064 24744
rect 19116 24692 19122 24744
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 21358 24732 21364 24744
rect 20027 24704 21364 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 21358 24692 21364 24704
rect 21416 24692 21422 24744
rect 22186 24664 22192 24676
rect 21008 24636 22192 24664
rect 21008 24596 21036 24636
rect 22186 24624 22192 24636
rect 22244 24624 22250 24676
rect 22480 24664 22508 24772
rect 22646 24692 22652 24744
rect 22704 24732 22710 24744
rect 22833 24735 22891 24741
rect 22833 24732 22845 24735
rect 22704 24704 22845 24732
rect 22704 24692 22710 24704
rect 22833 24701 22845 24704
rect 22879 24701 22891 24735
rect 22833 24695 22891 24701
rect 22925 24735 22983 24741
rect 22925 24701 22937 24735
rect 22971 24701 22983 24735
rect 22925 24695 22983 24701
rect 22940 24664 22968 24695
rect 23290 24692 23296 24744
rect 23348 24732 23354 24744
rect 23569 24735 23627 24741
rect 23569 24732 23581 24735
rect 23348 24704 23581 24732
rect 23348 24692 23354 24704
rect 23569 24701 23581 24704
rect 23615 24701 23627 24735
rect 23569 24695 23627 24701
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 23934 24732 23940 24744
rect 23891 24704 23940 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 23934 24692 23940 24704
rect 23992 24692 23998 24744
rect 22480 24636 22968 24664
rect 18984 24568 21036 24596
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 21453 24599 21511 24605
rect 21453 24596 21465 24599
rect 21324 24568 21465 24596
rect 21324 24556 21330 24568
rect 21453 24565 21465 24568
rect 21499 24565 21511 24599
rect 21453 24559 21511 24565
rect 22094 24556 22100 24608
rect 22152 24556 22158 24608
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 25222 24556 25228 24608
rect 25280 24596 25286 24608
rect 25317 24599 25375 24605
rect 25317 24596 25329 24599
rect 25280 24568 25329 24596
rect 25280 24556 25286 24568
rect 25317 24565 25329 24568
rect 25363 24565 25375 24599
rect 25317 24559 25375 24565
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 10042 24352 10048 24404
rect 10100 24352 10106 24404
rect 14642 24392 14648 24404
rect 10428 24364 14648 24392
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24188 5779 24191
rect 6454 24188 6460 24200
rect 5767 24160 6460 24188
rect 5767 24157 5779 24160
rect 5721 24151 5779 24157
rect 6454 24148 6460 24160
rect 6512 24148 6518 24200
rect 6825 24191 6883 24197
rect 6825 24157 6837 24191
rect 6871 24157 6883 24191
rect 6825 24151 6883 24157
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24188 7987 24191
rect 9582 24188 9588 24200
rect 7975 24160 9588 24188
rect 7975 24157 7987 24160
rect 7929 24151 7987 24157
rect 6840 24120 6868 24151
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10428 24197 10456 24364
rect 14642 24352 14648 24364
rect 14700 24352 14706 24404
rect 15289 24395 15347 24401
rect 15289 24361 15301 24395
rect 15335 24392 15347 24395
rect 15654 24392 15660 24404
rect 15335 24364 15660 24392
rect 15335 24361 15347 24364
rect 15289 24355 15347 24361
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 20254 24392 20260 24404
rect 15764 24364 20260 24392
rect 14458 24284 14464 24336
rect 14516 24324 14522 24336
rect 14921 24327 14979 24333
rect 14921 24324 14933 24327
rect 14516 24296 14933 24324
rect 14516 24284 14522 24296
rect 14921 24293 14933 24296
rect 14967 24293 14979 24327
rect 14921 24287 14979 24293
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24256 10747 24259
rect 10870 24256 10876 24268
rect 10735 24228 10876 24256
rect 10735 24225 10747 24228
rect 10689 24219 10747 24225
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11514 24216 11520 24268
rect 11572 24216 11578 24268
rect 15764 24256 15792 24364
rect 20254 24352 20260 24364
rect 20312 24352 20318 24404
rect 21542 24352 21548 24404
rect 21600 24352 21606 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 25225 24395 25283 24401
rect 25225 24392 25237 24395
rect 25188 24364 25237 24392
rect 25188 24352 25194 24364
rect 25225 24361 25237 24364
rect 25271 24361 25283 24395
rect 25225 24355 25283 24361
rect 17126 24284 17132 24336
rect 17184 24324 17190 24336
rect 19702 24324 19708 24336
rect 17184 24296 19708 24324
rect 17184 24284 17190 24296
rect 19702 24284 19708 24296
rect 19760 24284 19766 24336
rect 14476 24228 15792 24256
rect 10413 24191 10471 24197
rect 10413 24157 10425 24191
rect 10459 24157 10471 24191
rect 10413 24151 10471 24157
rect 11238 24148 11244 24200
rect 11296 24148 11302 24200
rect 12618 24148 12624 24200
rect 12676 24148 12682 24200
rect 13078 24148 13084 24200
rect 13136 24188 13142 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 13136 24160 14289 24188
rect 13136 24148 13142 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 8573 24123 8631 24129
rect 8573 24120 8585 24123
rect 6840 24092 8585 24120
rect 8573 24089 8585 24092
rect 8619 24089 8631 24123
rect 8573 24083 8631 24089
rect 9401 24123 9459 24129
rect 9401 24089 9413 24123
rect 9447 24120 9459 24123
rect 14476 24120 14504 24228
rect 17034 24216 17040 24268
rect 17092 24256 17098 24268
rect 18693 24259 18751 24265
rect 18693 24256 18705 24259
rect 17092 24228 18705 24256
rect 17092 24216 17098 24228
rect 18693 24225 18705 24228
rect 18739 24225 18751 24259
rect 18693 24219 18751 24225
rect 18874 24216 18880 24268
rect 18932 24256 18938 24268
rect 20073 24259 20131 24265
rect 18932 24228 20024 24256
rect 18932 24216 18938 24228
rect 15378 24148 15384 24200
rect 15436 24188 15442 24200
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 15436 24160 15485 24188
rect 15436 24148 15442 24160
rect 15473 24157 15485 24160
rect 15519 24188 15531 24191
rect 17494 24188 17500 24200
rect 15519 24160 17500 24188
rect 15519 24157 15531 24160
rect 15473 24151 15531 24157
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 18414 24148 18420 24200
rect 18472 24188 18478 24200
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 18472 24160 19809 24188
rect 18472 24148 18478 24160
rect 19797 24157 19809 24160
rect 19843 24157 19855 24191
rect 19996 24188 20024 24228
rect 20073 24225 20085 24259
rect 20119 24256 20131 24259
rect 20990 24256 20996 24268
rect 20119 24228 20996 24256
rect 20119 24225 20131 24228
rect 20073 24219 20131 24225
rect 20990 24216 20996 24228
rect 21048 24216 21054 24268
rect 19996 24160 20668 24188
rect 19797 24151 19855 24157
rect 9447 24092 11928 24120
rect 9447 24089 9459 24092
rect 9401 24083 9459 24089
rect 6365 24055 6423 24061
rect 6365 24021 6377 24055
rect 6411 24052 6423 24055
rect 6914 24052 6920 24064
rect 6411 24024 6920 24052
rect 6411 24021 6423 24024
rect 6365 24015 6423 24021
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 7466 24012 7472 24064
rect 7524 24012 7530 24064
rect 10502 24012 10508 24064
rect 10560 24012 10566 24064
rect 11900 24052 11928 24092
rect 12820 24092 14504 24120
rect 15933 24123 15991 24129
rect 12820 24052 12848 24092
rect 15933 24089 15945 24123
rect 15979 24120 15991 24123
rect 20438 24120 20444 24132
rect 15979 24092 20444 24120
rect 15979 24089 15991 24092
rect 15933 24083 15991 24089
rect 20438 24080 20444 24092
rect 20496 24080 20502 24132
rect 20640 24120 20668 24160
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 20901 24191 20959 24197
rect 20901 24188 20913 24191
rect 20772 24160 20913 24188
rect 20772 24148 20778 24160
rect 20901 24157 20913 24160
rect 20947 24188 20959 24191
rect 21634 24188 21640 24200
rect 20947 24160 21640 24188
rect 20947 24157 20959 24160
rect 20901 24151 20959 24157
rect 21634 24148 21640 24160
rect 21692 24148 21698 24200
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21968 24160 22017 24188
rect 21968 24148 21974 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 24578 24148 24584 24200
rect 24636 24148 24642 24200
rect 21266 24120 21272 24132
rect 20640 24092 21272 24120
rect 21266 24080 21272 24092
rect 21324 24080 21330 24132
rect 22278 24080 22284 24132
rect 22336 24080 22342 24132
rect 23658 24120 23664 24132
rect 23506 24092 23664 24120
rect 23658 24080 23664 24092
rect 23716 24120 23722 24132
rect 25314 24120 25320 24132
rect 23716 24092 25320 24120
rect 23716 24080 23722 24092
rect 25314 24080 25320 24092
rect 25372 24080 25378 24132
rect 11900 24024 12848 24052
rect 12989 24055 13047 24061
rect 12989 24021 13001 24055
rect 13035 24052 13047 24055
rect 13446 24052 13452 24064
rect 13035 24024 13452 24052
rect 13035 24021 13047 24024
rect 12989 24015 13047 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 13541 24055 13599 24061
rect 13541 24021 13553 24055
rect 13587 24052 13599 24055
rect 13722 24052 13728 24064
rect 13587 24024 13728 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 15657 24055 15715 24061
rect 15657 24052 15669 24055
rect 13964 24024 15669 24052
rect 13964 24012 13970 24024
rect 15657 24021 15669 24024
rect 15703 24052 15715 24055
rect 16666 24052 16672 24064
rect 15703 24024 16672 24052
rect 15703 24021 15715 24024
rect 15657 24015 15715 24021
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 17218 24012 17224 24064
rect 17276 24012 17282 24064
rect 18141 24055 18199 24061
rect 18141 24021 18153 24055
rect 18187 24052 18199 24055
rect 18414 24052 18420 24064
rect 18187 24024 18420 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 18506 24012 18512 24064
rect 18564 24012 18570 24064
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 18782 24052 18788 24064
rect 18647 24024 18788 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 18782 24012 18788 24024
rect 18840 24052 18846 24064
rect 19150 24052 19156 24064
rect 18840 24024 19156 24052
rect 18840 24012 18846 24024
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 20346 24052 20352 24064
rect 19944 24024 20352 24052
rect 19944 24012 19950 24024
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 23753 24055 23811 24061
rect 23753 24021 23765 24055
rect 23799 24052 23811 24055
rect 23842 24052 23848 24064
rect 23799 24024 23848 24052
rect 23799 24021 23811 24024
rect 23753 24015 23811 24021
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 24026 24012 24032 24064
rect 24084 24012 24090 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 6454 23808 6460 23860
rect 6512 23808 6518 23860
rect 9122 23808 9128 23860
rect 9180 23808 9186 23860
rect 9585 23851 9643 23857
rect 9585 23817 9597 23851
rect 9631 23848 9643 23851
rect 10042 23848 10048 23860
rect 9631 23820 10048 23848
rect 9631 23817 9643 23820
rect 9585 23811 9643 23817
rect 10042 23808 10048 23820
rect 10100 23808 10106 23860
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 11149 23851 11207 23857
rect 11149 23848 11161 23851
rect 10376 23820 11161 23848
rect 10376 23808 10382 23820
rect 11149 23817 11161 23820
rect 11195 23817 11207 23851
rect 11149 23811 11207 23817
rect 11793 23851 11851 23857
rect 11793 23817 11805 23851
rect 11839 23817 11851 23851
rect 11793 23811 11851 23817
rect 6472 23576 6500 23808
rect 7650 23740 7656 23792
rect 7708 23780 7714 23792
rect 11808 23780 11836 23811
rect 13078 23808 13084 23860
rect 13136 23808 13142 23860
rect 13906 23808 13912 23860
rect 13964 23808 13970 23860
rect 15841 23851 15899 23857
rect 15841 23817 15853 23851
rect 15887 23848 15899 23851
rect 16022 23848 16028 23860
rect 15887 23820 16028 23848
rect 15887 23817 15899 23820
rect 15841 23811 15899 23817
rect 16022 23808 16028 23820
rect 16080 23808 16086 23860
rect 18506 23808 18512 23860
rect 18564 23848 18570 23860
rect 19242 23848 19248 23860
rect 18564 23820 19248 23848
rect 18564 23808 18570 23820
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 19518 23848 19524 23860
rect 19352 23820 19524 23848
rect 7708 23752 11836 23780
rect 7708 23740 7714 23752
rect 12066 23740 12072 23792
rect 12124 23780 12130 23792
rect 12124 23752 13952 23780
rect 12124 23740 12130 23752
rect 6914 23672 6920 23724
rect 6972 23672 6978 23724
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23712 9551 23715
rect 10318 23712 10324 23724
rect 9539 23684 10324 23712
rect 9539 23681 9551 23684
rect 9493 23675 9551 23681
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 11977 23715 12035 23721
rect 11977 23681 11989 23715
rect 12023 23681 12035 23715
rect 11977 23675 12035 23681
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 13924 23712 13952 23752
rect 13998 23740 14004 23792
rect 14056 23740 14062 23792
rect 19352 23789 19380 23820
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19702 23808 19708 23860
rect 19760 23848 19766 23860
rect 21821 23851 21879 23857
rect 21821 23848 21833 23851
rect 19760 23820 21833 23848
rect 19760 23808 19766 23820
rect 21821 23817 21833 23820
rect 21867 23848 21879 23851
rect 22373 23851 22431 23857
rect 22373 23848 22385 23851
rect 21867 23820 22385 23848
rect 21867 23817 21879 23820
rect 21821 23811 21879 23817
rect 22373 23817 22385 23820
rect 22419 23817 22431 23851
rect 22373 23811 22431 23817
rect 22465 23851 22523 23857
rect 22465 23817 22477 23851
rect 22511 23848 22523 23851
rect 24210 23848 24216 23860
rect 22511 23820 24216 23848
rect 22511 23817 22523 23820
rect 22465 23811 22523 23817
rect 24210 23808 24216 23820
rect 24268 23808 24274 23860
rect 24946 23808 24952 23860
rect 25004 23848 25010 23860
rect 25406 23848 25412 23860
rect 25004 23820 25412 23848
rect 25004 23808 25010 23820
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 19337 23783 19395 23789
rect 19337 23749 19349 23783
rect 19383 23749 19395 23783
rect 23382 23780 23388 23792
rect 20562 23752 21864 23780
rect 19337 23743 19395 23749
rect 12483 23684 13860 23712
rect 13924 23684 14228 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 7190 23604 7196 23656
rect 7248 23604 7254 23656
rect 9674 23604 9680 23656
rect 9732 23604 9738 23656
rect 10134 23604 10140 23656
rect 10192 23644 10198 23656
rect 10520 23644 10548 23675
rect 10192 23616 10548 23644
rect 11992 23644 12020 23675
rect 12802 23644 12808 23656
rect 11992 23616 12808 23644
rect 10192 23604 10198 23616
rect 12802 23604 12808 23616
rect 12860 23604 12866 23656
rect 13262 23576 13268 23588
rect 6472 23548 13268 23576
rect 13262 23536 13268 23548
rect 13320 23536 13326 23588
rect 8297 23511 8355 23517
rect 8297 23477 8309 23511
rect 8343 23508 8355 23511
rect 8386 23508 8392 23520
rect 8343 23480 8392 23508
rect 8343 23477 8355 23480
rect 8297 23471 8355 23477
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 12618 23468 12624 23520
rect 12676 23508 12682 23520
rect 13541 23511 13599 23517
rect 13541 23508 13553 23511
rect 12676 23480 13553 23508
rect 12676 23468 12682 23480
rect 13541 23477 13553 23480
rect 13587 23477 13599 23511
rect 13832 23508 13860 23684
rect 14200 23653 14228 23684
rect 14642 23672 14648 23724
rect 14700 23712 14706 23724
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 14700 23684 14749 23712
rect 14700 23672 14706 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 17957 23715 18015 23721
rect 17957 23681 17969 23715
rect 18003 23712 18015 23715
rect 18003 23684 19012 23712
rect 18003 23681 18015 23684
rect 17957 23675 18015 23681
rect 14185 23647 14243 23653
rect 14185 23613 14197 23647
rect 14231 23613 14243 23647
rect 18984 23644 19012 23684
rect 19058 23672 19064 23724
rect 19116 23672 19122 23724
rect 20070 23644 20076 23656
rect 18984 23616 20076 23644
rect 14185 23607 14243 23613
rect 20070 23604 20076 23616
rect 20128 23644 20134 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20128 23616 20821 23644
rect 20128 23604 20134 23616
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 20809 23607 20867 23613
rect 21100 23520 21128 23752
rect 21836 23724 21864 23752
rect 23124 23752 23388 23780
rect 21450 23672 21456 23724
rect 21508 23672 21514 23724
rect 21818 23672 21824 23724
rect 21876 23672 21882 23724
rect 22646 23604 22652 23656
rect 22704 23644 22710 23656
rect 23124 23644 23152 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 25314 23780 25320 23792
rect 24702 23752 25320 23780
rect 25314 23740 25320 23752
rect 25372 23780 25378 23792
rect 25501 23783 25559 23789
rect 25501 23780 25513 23783
rect 25372 23752 25513 23780
rect 25372 23740 25378 23752
rect 25501 23749 25513 23752
rect 25547 23749 25559 23783
rect 25501 23743 25559 23749
rect 22704 23616 23152 23644
rect 22704 23604 22710 23616
rect 23198 23604 23204 23656
rect 23256 23604 23262 23656
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 25682 23644 25688 23656
rect 23523 23616 25688 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 25682 23604 25688 23616
rect 25740 23604 25746 23656
rect 21450 23536 21456 23588
rect 21508 23576 21514 23588
rect 21910 23576 21916 23588
rect 21508 23548 21916 23576
rect 21508 23536 21514 23548
rect 21910 23536 21916 23548
rect 21968 23576 21974 23588
rect 23216 23576 23244 23604
rect 21968 23548 23244 23576
rect 21968 23536 21974 23548
rect 15381 23511 15439 23517
rect 15381 23508 15393 23511
rect 13832 23480 15393 23508
rect 13541 23471 13599 23477
rect 15381 23477 15393 23480
rect 15427 23477 15439 23511
rect 15381 23471 15439 23477
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 17497 23511 17555 23517
rect 17497 23508 17509 23511
rect 15528 23480 17509 23508
rect 15528 23468 15534 23480
rect 17497 23477 17509 23480
rect 17543 23477 17555 23511
rect 17497 23471 17555 23477
rect 18601 23511 18659 23517
rect 18601 23477 18613 23511
rect 18647 23508 18659 23511
rect 20622 23508 20628 23520
rect 18647 23480 20628 23508
rect 18647 23477 18659 23480
rect 18601 23471 18659 23477
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 21082 23468 21088 23520
rect 21140 23468 21146 23520
rect 21266 23468 21272 23520
rect 21324 23468 21330 23520
rect 22002 23468 22008 23520
rect 22060 23468 22066 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 8478 23264 8484 23316
rect 8536 23304 8542 23316
rect 8573 23307 8631 23313
rect 8573 23304 8585 23307
rect 8536 23276 8585 23304
rect 8536 23264 8542 23276
rect 8573 23273 8585 23276
rect 8619 23273 8631 23307
rect 8573 23267 8631 23273
rect 9232 23276 10456 23304
rect 7193 23239 7251 23245
rect 7193 23205 7205 23239
rect 7239 23236 7251 23239
rect 9232 23236 9260 23276
rect 7239 23208 9260 23236
rect 10428 23236 10456 23276
rect 12802 23264 12808 23316
rect 12860 23304 12866 23316
rect 12989 23307 13047 23313
rect 12989 23304 13001 23307
rect 12860 23276 13001 23304
rect 12860 23264 12866 23276
rect 12989 23273 13001 23276
rect 13035 23273 13047 23307
rect 21542 23304 21548 23316
rect 12989 23267 13047 23273
rect 14384 23276 21548 23304
rect 14384 23236 14412 23276
rect 21542 23264 21548 23276
rect 21600 23264 21606 23316
rect 21818 23264 21824 23316
rect 21876 23304 21882 23316
rect 22281 23307 22339 23313
rect 22281 23304 22293 23307
rect 21876 23276 22293 23304
rect 21876 23264 21882 23276
rect 22281 23273 22293 23276
rect 22327 23304 22339 23307
rect 23658 23304 23664 23316
rect 22327 23276 23664 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 23658 23264 23664 23276
rect 23716 23264 23722 23316
rect 10428 23208 14412 23236
rect 7239 23205 7251 23208
rect 7193 23199 7251 23205
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23168 6055 23171
rect 7650 23168 7656 23180
rect 6043 23140 7656 23168
rect 6043 23137 6055 23140
rect 5997 23131 6055 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 6270 23060 6276 23112
rect 6328 23060 6334 23112
rect 7285 23103 7343 23109
rect 7285 23069 7297 23103
rect 7331 23100 7343 23103
rect 7760 23100 7788 23208
rect 16482 23196 16488 23248
rect 16540 23236 16546 23248
rect 18877 23239 18935 23245
rect 16540 23208 17172 23236
rect 16540 23196 16546 23208
rect 7834 23128 7840 23180
rect 7892 23168 7898 23180
rect 9125 23171 9183 23177
rect 9125 23168 9137 23171
rect 7892 23140 9137 23168
rect 7892 23128 7898 23140
rect 9125 23137 9137 23140
rect 9171 23137 9183 23171
rect 9125 23131 9183 23137
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 9456 23140 10640 23168
rect 9456 23128 9462 23140
rect 7331 23072 7788 23100
rect 7929 23103 7987 23109
rect 7331 23069 7343 23072
rect 7285 23063 7343 23069
rect 7929 23069 7941 23103
rect 7975 23069 7987 23103
rect 10612 23100 10640 23140
rect 10686 23128 10692 23180
rect 10744 23168 10750 23180
rect 12253 23171 12311 23177
rect 12253 23168 12265 23171
rect 10744 23140 12265 23168
rect 10744 23128 10750 23140
rect 12253 23137 12265 23140
rect 12299 23137 12311 23171
rect 12253 23131 12311 23137
rect 13446 23128 13452 23180
rect 13504 23168 13510 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13504 23140 13553 23168
rect 13504 23128 13510 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 13541 23131 13599 23137
rect 14553 23171 14611 23177
rect 14553 23137 14565 23171
rect 14599 23168 14611 23171
rect 15194 23168 15200 23180
rect 14599 23140 15200 23168
rect 14599 23137 14611 23140
rect 14553 23131 14611 23137
rect 15194 23128 15200 23140
rect 15252 23128 15258 23180
rect 15930 23128 15936 23180
rect 15988 23168 15994 23180
rect 17037 23171 17095 23177
rect 17037 23168 17049 23171
rect 15988 23140 17049 23168
rect 15988 23128 15994 23140
rect 17037 23137 17049 23140
rect 17083 23137 17095 23171
rect 17037 23131 17095 23137
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 10612 23072 12081 23100
rect 7929 23063 7987 23069
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23100 12219 23103
rect 12526 23100 12532 23112
rect 12207 23072 12532 23100
rect 12207 23069 12219 23072
rect 12161 23063 12219 23069
rect 7944 22964 7972 23063
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 12636 23072 13492 23100
rect 9401 23035 9459 23041
rect 9401 23001 9413 23035
rect 9447 23032 9459 23035
rect 9674 23032 9680 23044
rect 9447 23004 9680 23032
rect 9447 23001 9459 23004
rect 9401 22995 9459 23001
rect 9674 22992 9680 23004
rect 9732 22992 9738 23044
rect 10778 23032 10784 23044
rect 10626 23004 10784 23032
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 12636 23032 12664 23072
rect 13357 23035 13415 23041
rect 13357 23032 13369 23035
rect 11716 23004 12664 23032
rect 12728 23004 13369 23032
rect 10870 22964 10876 22976
rect 7944 22936 10876 22964
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 11716 22973 11744 23004
rect 11701 22967 11759 22973
rect 11701 22933 11713 22967
rect 11747 22933 11759 22967
rect 11701 22927 11759 22933
rect 12158 22924 12164 22976
rect 12216 22964 12222 22976
rect 12728 22964 12756 23004
rect 13357 23001 13369 23004
rect 13403 23001 13415 23035
rect 13464 23032 13492 23072
rect 14274 23060 14280 23112
rect 14332 23060 14338 23112
rect 16945 23103 17003 23109
rect 16945 23069 16957 23103
rect 16991 23100 17003 23103
rect 17144 23100 17172 23208
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 21634 23236 21640 23248
rect 18923 23208 21640 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 21634 23196 21640 23208
rect 21692 23196 21698 23248
rect 17773 23171 17831 23177
rect 17773 23137 17785 23171
rect 17819 23168 17831 23171
rect 18598 23168 18604 23180
rect 17819 23140 18604 23168
rect 17819 23137 17831 23140
rect 17773 23131 17831 23137
rect 17788 23100 17816 23131
rect 18598 23128 18604 23140
rect 18656 23128 18662 23180
rect 19334 23128 19340 23180
rect 19392 23128 19398 23180
rect 19610 23128 19616 23180
rect 19668 23168 19674 23180
rect 19886 23168 19892 23180
rect 19668 23140 19892 23168
rect 19668 23128 19674 23140
rect 19886 23128 19892 23140
rect 19944 23128 19950 23180
rect 20533 23171 20591 23177
rect 20533 23137 20545 23171
rect 20579 23168 20591 23171
rect 20714 23168 20720 23180
rect 20579 23140 20720 23168
rect 20579 23137 20591 23140
rect 20533 23131 20591 23137
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 22097 23171 22155 23177
rect 22097 23168 22109 23171
rect 20864 23140 22109 23168
rect 20864 23128 20870 23140
rect 22097 23137 22109 23140
rect 22143 23137 22155 23171
rect 22097 23131 22155 23137
rect 23845 23171 23903 23177
rect 23845 23137 23857 23171
rect 23891 23168 23903 23171
rect 24486 23168 24492 23180
rect 23891 23140 24492 23168
rect 23891 23137 23903 23140
rect 23845 23131 23903 23137
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 16991 23072 17816 23100
rect 18233 23103 18291 23109
rect 16991 23069 17003 23072
rect 16945 23063 17003 23069
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 20162 23100 20168 23112
rect 18279 23072 20168 23100
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 20162 23060 20168 23072
rect 20220 23060 20226 23112
rect 20254 23060 20260 23112
rect 20312 23060 20318 23112
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 21085 23103 21143 23109
rect 21085 23100 21097 23103
rect 20680 23072 21097 23100
rect 20680 23060 20686 23072
rect 21085 23069 21097 23072
rect 21131 23069 21143 23103
rect 21085 23063 21143 23069
rect 21818 23060 21824 23112
rect 21876 23100 21882 23112
rect 22649 23103 22707 23109
rect 22649 23100 22661 23103
rect 21876 23072 22661 23100
rect 21876 23060 21882 23072
rect 22649 23069 22661 23072
rect 22695 23069 22707 23103
rect 22649 23063 22707 23069
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23100 25099 23103
rect 25590 23100 25596 23112
rect 25087 23072 25596 23100
rect 25087 23069 25099 23072
rect 25041 23063 25099 23069
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 13464 23004 14964 23032
rect 13357 22995 13415 23001
rect 12216 22936 12756 22964
rect 13449 22967 13507 22973
rect 12216 22924 12222 22936
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 14734 22964 14740 22976
rect 13495 22936 14740 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 14936 22964 14964 23004
rect 15010 22992 15016 23044
rect 15068 22992 15074 23044
rect 20349 23035 20407 23041
rect 20349 23001 20361 23035
rect 20395 23032 20407 23035
rect 23382 23032 23388 23044
rect 20395 23004 23388 23032
rect 20395 23001 20407 23004
rect 20349 22995 20407 23001
rect 23382 22992 23388 23004
rect 23440 22992 23446 23044
rect 24949 23035 25007 23041
rect 24949 23001 24961 23035
rect 24995 23032 25007 23035
rect 25774 23032 25780 23044
rect 24995 23004 25780 23032
rect 24995 23001 25007 23004
rect 24949 22995 25007 23001
rect 25774 22992 25780 23004
rect 25832 23032 25838 23044
rect 26142 23032 26148 23044
rect 25832 23004 26148 23032
rect 25832 22992 25838 23004
rect 26142 22992 26148 23004
rect 26200 22992 26206 23044
rect 15838 22964 15844 22976
rect 14936 22936 15844 22964
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16025 22967 16083 22973
rect 16025 22933 16037 22967
rect 16071 22964 16083 22967
rect 16114 22964 16120 22976
rect 16071 22936 16120 22964
rect 16071 22933 16083 22936
rect 16025 22927 16083 22933
rect 16114 22924 16120 22936
rect 16172 22924 16178 22976
rect 16482 22924 16488 22976
rect 16540 22924 16546 22976
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 16853 22967 16911 22973
rect 16853 22964 16865 22967
rect 16724 22936 16865 22964
rect 16724 22924 16730 22936
rect 16853 22933 16865 22936
rect 16899 22964 16911 22967
rect 17589 22967 17647 22973
rect 17589 22964 17601 22967
rect 16899 22936 17601 22964
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 17589 22933 17601 22936
rect 17635 22964 17647 22967
rect 17862 22964 17868 22976
rect 17635 22936 17868 22964
rect 17635 22933 17647 22936
rect 17589 22927 17647 22933
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 17957 22967 18015 22973
rect 17957 22933 17969 22967
rect 18003 22964 18015 22967
rect 18782 22964 18788 22976
rect 18003 22936 18788 22964
rect 18003 22933 18015 22936
rect 17957 22927 18015 22933
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 19521 22967 19579 22973
rect 19521 22933 19533 22967
rect 19567 22964 19579 22967
rect 19610 22964 19616 22976
rect 19567 22936 19616 22964
rect 19567 22933 19579 22936
rect 19521 22927 19579 22933
rect 19610 22924 19616 22936
rect 19668 22924 19674 22976
rect 19886 22924 19892 22976
rect 19944 22924 19950 22976
rect 20714 22924 20720 22976
rect 20772 22964 20778 22976
rect 21729 22967 21787 22973
rect 21729 22964 21741 22967
rect 20772 22936 21741 22964
rect 20772 22924 20778 22936
rect 21729 22933 21741 22936
rect 21775 22933 21787 22967
rect 21729 22927 21787 22933
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22964 24639 22967
rect 24670 22964 24676 22976
rect 24627 22936 24676 22964
rect 24627 22933 24639 22936
rect 24581 22927 24639 22933
rect 24670 22924 24676 22936
rect 24728 22924 24734 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 12069 22763 12127 22769
rect 12069 22729 12081 22763
rect 12115 22760 12127 22763
rect 12342 22760 12348 22772
rect 12115 22732 12348 22760
rect 12115 22729 12127 22732
rect 12069 22723 12127 22729
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 14918 22760 14924 22772
rect 14016 22732 14924 22760
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22692 6699 22695
rect 9122 22692 9128 22704
rect 6687 22664 9128 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 10134 22692 10140 22704
rect 10074 22664 10140 22692
rect 10134 22652 10140 22664
rect 10192 22692 10198 22704
rect 10778 22692 10784 22704
rect 10192 22664 10784 22692
rect 10192 22652 10198 22664
rect 10778 22652 10784 22664
rect 10836 22652 10842 22704
rect 12161 22695 12219 22701
rect 12161 22661 12173 22695
rect 12207 22692 12219 22695
rect 13354 22692 13360 22704
rect 12207 22664 13360 22692
rect 12207 22661 12219 22664
rect 12161 22655 12219 22661
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7834 22624 7840 22636
rect 7248 22596 7840 22624
rect 7248 22584 7254 22596
rect 7834 22584 7840 22596
rect 7892 22624 7898 22636
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 7892 22596 8585 22624
rect 7892 22584 7898 22596
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 12897 22627 12955 22633
rect 12897 22593 12909 22627
rect 12943 22624 12955 22627
rect 14016 22624 14044 22732
rect 14918 22720 14924 22732
rect 14976 22760 14982 22772
rect 15749 22763 15807 22769
rect 15749 22760 15761 22763
rect 14976 22732 15761 22760
rect 14976 22720 14982 22732
rect 15749 22729 15761 22732
rect 15795 22760 15807 22763
rect 16206 22760 16212 22772
rect 15795 22732 16212 22760
rect 15795 22729 15807 22732
rect 15749 22723 15807 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 16850 22720 16856 22772
rect 16908 22760 16914 22772
rect 17497 22763 17555 22769
rect 17497 22760 17509 22763
rect 16908 22732 17509 22760
rect 16908 22720 16914 22732
rect 17497 22729 17509 22732
rect 17543 22729 17555 22763
rect 17497 22723 17555 22729
rect 18417 22763 18475 22769
rect 18417 22729 18429 22763
rect 18463 22760 18475 22763
rect 18690 22760 18696 22772
rect 18463 22732 18696 22760
rect 18463 22729 18475 22732
rect 18417 22723 18475 22729
rect 18690 22720 18696 22732
rect 18748 22760 18754 22772
rect 19150 22760 19156 22772
rect 18748 22732 19156 22760
rect 18748 22720 18754 22732
rect 19150 22720 19156 22732
rect 19208 22720 19214 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 19889 22763 19947 22769
rect 19889 22760 19901 22763
rect 19484 22732 19901 22760
rect 19484 22720 19490 22732
rect 19889 22729 19901 22732
rect 19935 22729 19947 22763
rect 19889 22723 19947 22729
rect 19981 22763 20039 22769
rect 19981 22729 19993 22763
rect 20027 22760 20039 22763
rect 20898 22760 20904 22772
rect 20027 22732 20904 22760
rect 20027 22729 20039 22732
rect 19981 22723 20039 22729
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 21358 22720 21364 22772
rect 21416 22720 21422 22772
rect 14734 22652 14740 22704
rect 14792 22652 14798 22704
rect 15838 22652 15844 22704
rect 15896 22692 15902 22704
rect 18230 22692 18236 22704
rect 15896 22664 18236 22692
rect 15896 22652 15902 22664
rect 18230 22652 18236 22664
rect 18288 22652 18294 22704
rect 18322 22652 18328 22704
rect 18380 22692 18386 22704
rect 18969 22695 19027 22701
rect 18969 22692 18981 22695
rect 18380 22664 18981 22692
rect 18380 22652 18386 22664
rect 18969 22661 18981 22664
rect 19015 22692 19027 22695
rect 19058 22692 19064 22704
rect 19015 22664 19064 22692
rect 19015 22661 19027 22664
rect 18969 22655 19027 22661
rect 19058 22652 19064 22664
rect 19116 22652 19122 22704
rect 21726 22652 21732 22704
rect 21784 22692 21790 22704
rect 21784 22664 23980 22692
rect 21784 22652 21790 22664
rect 12943 22596 14044 22624
rect 12943 22593 12955 22596
rect 12897 22587 12955 22593
rect 16666 22584 16672 22636
rect 16724 22624 16730 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16724 22596 16865 22624
rect 16724 22584 16730 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 20714 22584 20720 22636
rect 20772 22584 20778 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 23952 22633 23980 22664
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 24946 22624 24952 22636
rect 23937 22587 23995 22593
rect 24688 22596 24952 22624
rect 7285 22559 7343 22565
rect 7285 22525 7297 22559
rect 7331 22525 7343 22559
rect 7285 22519 7343 22525
rect 7561 22559 7619 22565
rect 7561 22525 7573 22559
rect 7607 22556 7619 22559
rect 7650 22556 7656 22568
rect 7607 22528 7656 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 7193 22491 7251 22497
rect 7193 22457 7205 22491
rect 7239 22488 7251 22491
rect 7300 22488 7328 22519
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 8846 22516 8852 22568
rect 8904 22516 8910 22568
rect 10962 22516 10968 22568
rect 11020 22516 11026 22568
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22525 12311 22559
rect 12253 22519 12311 22525
rect 14001 22559 14059 22565
rect 14001 22525 14013 22559
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 14277 22559 14335 22565
rect 14277 22525 14289 22559
rect 14323 22556 14335 22559
rect 15470 22556 15476 22568
rect 14323 22528 15476 22556
rect 14323 22525 14335 22528
rect 14277 22519 14335 22525
rect 8478 22488 8484 22500
rect 7239 22460 8484 22488
rect 7239 22457 7251 22460
rect 7193 22451 7251 22457
rect 8478 22448 8484 22460
rect 8536 22448 8542 22500
rect 12268 22488 12296 22519
rect 10336 22460 12296 22488
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 10336 22429 10364 22460
rect 10321 22423 10379 22429
rect 10321 22420 10333 22423
rect 7892 22392 10333 22420
rect 7892 22380 7898 22392
rect 10321 22389 10333 22392
rect 10367 22389 10379 22423
rect 10321 22383 10379 22389
rect 10686 22380 10692 22432
rect 10744 22380 10750 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11112 22392 11713 22420
rect 11112 22380 11118 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 13538 22380 13544 22432
rect 13596 22380 13602 22432
rect 14016 22420 14044 22519
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 16390 22516 16396 22568
rect 16448 22516 16454 22568
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 18509 22559 18567 22565
rect 18509 22556 18521 22559
rect 17552 22528 18521 22556
rect 17552 22516 17558 22528
rect 18509 22525 18521 22528
rect 18555 22525 18567 22559
rect 18509 22519 18567 22525
rect 20070 22516 20076 22568
rect 20128 22516 20134 22568
rect 23293 22559 23351 22565
rect 23293 22525 23305 22559
rect 23339 22556 23351 22559
rect 24688 22556 24716 22596
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 23339 22528 24716 22556
rect 23339 22525 23351 22528
rect 23293 22519 23351 22525
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 16850 22488 16856 22500
rect 15304 22460 16856 22488
rect 14274 22420 14280 22432
rect 14016 22392 14280 22420
rect 14274 22380 14280 22392
rect 14332 22420 14338 22432
rect 15304 22420 15332 22460
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 20162 22448 20168 22500
rect 20220 22488 20226 22500
rect 26050 22488 26056 22500
rect 20220 22460 26056 22488
rect 20220 22448 20226 22460
rect 26050 22448 26056 22460
rect 26108 22448 26114 22500
rect 14332 22392 15332 22420
rect 17957 22423 18015 22429
rect 14332 22380 14338 22392
rect 17957 22389 17969 22423
rect 18003 22420 18015 22423
rect 18690 22420 18696 22432
rect 18003 22392 18696 22420
rect 18003 22389 18015 22392
rect 17957 22383 18015 22389
rect 18690 22380 18696 22392
rect 18748 22380 18754 22432
rect 19518 22380 19524 22432
rect 19576 22380 19582 22432
rect 25314 22380 25320 22432
rect 25372 22420 25378 22432
rect 25590 22420 25596 22432
rect 25372 22392 25596 22420
rect 25372 22380 25378 22392
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 6270 22176 6276 22228
rect 6328 22216 6334 22228
rect 15102 22216 15108 22228
rect 6328 22188 15108 22216
rect 6328 22176 6334 22188
rect 15102 22176 15108 22188
rect 15160 22176 15166 22228
rect 19242 22176 19248 22228
rect 19300 22176 19306 22228
rect 20162 22176 20168 22228
rect 20220 22216 20226 22228
rect 20993 22219 21051 22225
rect 20993 22216 21005 22219
rect 20220 22188 21005 22216
rect 20220 22176 20226 22188
rect 20993 22185 21005 22188
rect 21039 22216 21051 22219
rect 21082 22216 21088 22228
rect 21039 22188 21088 22216
rect 21039 22185 21051 22188
rect 20993 22179 21051 22185
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 21716 22219 21774 22225
rect 21716 22185 21728 22219
rect 21762 22216 21774 22219
rect 25314 22216 25320 22228
rect 21762 22188 25320 22216
rect 21762 22185 21774 22188
rect 21716 22179 21774 22185
rect 25314 22176 25320 22188
rect 25372 22176 25378 22228
rect 10594 22108 10600 22160
rect 10652 22148 10658 22160
rect 10652 22120 10824 22148
rect 10652 22108 10658 22120
rect 10796 22094 10824 22120
rect 13354 22108 13360 22160
rect 13412 22148 13418 22160
rect 13412 22120 15332 22148
rect 13412 22108 13418 22120
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22080 6883 22083
rect 7098 22080 7104 22092
rect 6871 22052 7104 22080
rect 6871 22049 6883 22052
rect 6825 22043 6883 22049
rect 7098 22040 7104 22052
rect 7156 22040 7162 22092
rect 10796 22089 10861 22094
rect 8573 22083 8631 22089
rect 8573 22049 8585 22083
rect 8619 22049 8631 22083
rect 8573 22043 8631 22049
rect 10781 22083 10861 22089
rect 10781 22049 10793 22083
rect 10827 22066 10861 22083
rect 13446 22080 13452 22092
rect 10827 22049 10839 22066
rect 10781 22043 10839 22049
rect 12406 22052 13452 22080
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 6181 21879 6239 21885
rect 6181 21876 6193 21879
rect 3752 21848 6193 21876
rect 3752 21836 3758 21848
rect 6181 21845 6193 21848
rect 6227 21845 6239 21879
rect 6380 21876 6408 21975
rect 8202 21972 8208 22024
rect 8260 21972 8266 22024
rect 8588 22012 8616 22043
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8588 21984 9137 22012
rect 9125 21981 9137 21984
rect 9171 22012 9183 22015
rect 9582 22012 9588 22024
rect 9171 21984 9588 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10686 22012 10692 22024
rect 10008 21984 10692 22012
rect 10008 21972 10014 21984
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 22012 12035 22015
rect 12406 22012 12434 22052
rect 13446 22040 13452 22052
rect 13504 22040 13510 22092
rect 13814 22040 13820 22092
rect 13872 22080 13878 22092
rect 15304 22089 15332 22120
rect 15289 22083 15347 22089
rect 13872 22052 15240 22080
rect 13872 22040 13878 22052
rect 12023 21984 12434 22012
rect 13081 22015 13139 22021
rect 12023 21981 12035 21984
rect 11977 21975 12035 21981
rect 13081 21981 13093 22015
rect 13127 22012 13139 22015
rect 13538 22012 13544 22024
rect 13127 21984 13544 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 13538 21972 13544 21984
rect 13596 21972 13602 22024
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 13780 21984 15117 22012
rect 13780 21972 13786 21984
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 15212 22012 15240 22052
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 16485 22083 16543 22089
rect 16485 22080 16497 22083
rect 16172 22052 16497 22080
rect 16172 22040 16178 22052
rect 16485 22049 16497 22052
rect 16531 22049 16543 22083
rect 16485 22043 16543 22049
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 15212 21984 16313 22012
rect 15105 21975 15163 21981
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 16574 22012 16580 22024
rect 16439 21984 16580 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 17494 22012 17500 22024
rect 17175 21984 17500 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 22012 18291 22015
rect 18782 22012 18788 22024
rect 18279 21984 18788 22012
rect 18279 21981 18291 21984
rect 18233 21975 18291 21981
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 19260 22012 19288 22176
rect 19334 22040 19340 22092
rect 19392 22080 19398 22092
rect 19429 22083 19487 22089
rect 19429 22080 19441 22083
rect 19392 22052 19441 22080
rect 19392 22040 19398 22052
rect 19429 22049 19441 22052
rect 19475 22080 19487 22083
rect 20441 22083 20499 22089
rect 19475 22052 20208 22080
rect 19475 22049 19487 22052
rect 19429 22043 19487 22049
rect 20180 22021 20208 22052
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 20487 22052 20944 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 20165 22015 20223 22021
rect 19260 21984 19380 22012
rect 6730 21904 6736 21956
rect 6788 21944 6794 21956
rect 7101 21947 7159 21953
rect 7101 21944 7113 21947
rect 6788 21916 7113 21944
rect 6788 21904 6794 21916
rect 7101 21913 7113 21916
rect 7147 21913 7159 21947
rect 7101 21907 7159 21913
rect 8496 21916 15976 21944
rect 8496 21876 8524 21916
rect 6380 21848 8524 21876
rect 6181 21839 6239 21845
rect 8662 21836 8668 21888
rect 8720 21876 8726 21888
rect 9769 21879 9827 21885
rect 9769 21876 9781 21879
rect 8720 21848 9781 21876
rect 8720 21836 8726 21848
rect 9769 21845 9781 21848
rect 9815 21845 9827 21879
rect 9769 21839 9827 21845
rect 10226 21836 10232 21888
rect 10284 21836 10290 21888
rect 10594 21836 10600 21888
rect 10652 21836 10658 21888
rect 10778 21836 10784 21888
rect 10836 21876 10842 21888
rect 11517 21879 11575 21885
rect 11517 21876 11529 21879
rect 10836 21848 11529 21876
rect 10836 21836 10842 21848
rect 11517 21845 11529 21848
rect 11563 21845 11575 21879
rect 11517 21839 11575 21845
rect 12618 21836 12624 21888
rect 12676 21836 12682 21888
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 13725 21879 13783 21885
rect 13725 21876 13737 21879
rect 13228 21848 13737 21876
rect 13228 21836 13234 21848
rect 13725 21845 13737 21848
rect 13771 21845 13783 21879
rect 13725 21839 13783 21845
rect 14550 21836 14556 21888
rect 14608 21876 14614 21888
rect 14737 21879 14795 21885
rect 14737 21876 14749 21879
rect 14608 21848 14749 21876
rect 14608 21836 14614 21848
rect 14737 21845 14749 21848
rect 14783 21845 14795 21879
rect 14737 21839 14795 21845
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 15948 21885 15976 21916
rect 17862 21904 17868 21956
rect 17920 21944 17926 21956
rect 19242 21944 19248 21956
rect 17920 21916 19248 21944
rect 17920 21904 17926 21916
rect 19242 21904 19248 21916
rect 19300 21904 19306 21956
rect 19352 21944 19380 21984
rect 20165 21981 20177 22015
rect 20211 21981 20223 22015
rect 20165 21975 20223 21981
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 22012 20315 22015
rect 20806 22012 20812 22024
rect 20303 21984 20812 22012
rect 20303 21981 20315 21984
rect 20257 21975 20315 21981
rect 20272 21944 20300 21975
rect 20806 21972 20812 21984
rect 20864 21972 20870 22024
rect 19352 21916 20300 21944
rect 15197 21879 15255 21885
rect 15197 21876 15209 21879
rect 15160 21848 15209 21876
rect 15160 21836 15166 21848
rect 15197 21845 15209 21848
rect 15243 21845 15255 21879
rect 15197 21839 15255 21845
rect 15933 21879 15991 21885
rect 15933 21845 15945 21879
rect 15979 21845 15991 21879
rect 15933 21839 15991 21845
rect 17770 21836 17776 21888
rect 17828 21836 17834 21888
rect 18874 21836 18880 21888
rect 18932 21836 18938 21888
rect 19797 21879 19855 21885
rect 19797 21845 19809 21879
rect 19843 21876 19855 21879
rect 20806 21876 20812 21888
rect 19843 21848 20812 21876
rect 19843 21845 19855 21848
rect 19797 21839 19855 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 20916 21876 20944 22052
rect 21450 22040 21456 22092
rect 21508 22040 21514 22092
rect 21726 22040 21732 22092
rect 21784 22080 21790 22092
rect 21784 22052 23980 22080
rect 21784 22040 21790 22052
rect 21082 21972 21088 22024
rect 21140 21972 21146 22024
rect 23952 22021 23980 22052
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 24486 22080 24492 22092
rect 24084 22052 24492 22080
rect 24084 22040 24090 22052
rect 24486 22040 24492 22052
rect 24544 22040 24550 22092
rect 25038 22040 25044 22092
rect 25096 22040 25102 22092
rect 25222 22040 25228 22092
rect 25280 22040 25286 22092
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 21100 21944 21128 21972
rect 22002 21944 22008 21956
rect 21100 21916 22008 21944
rect 22002 21904 22008 21916
rect 22060 21944 22066 21956
rect 22060 21916 22218 21944
rect 22060 21904 22066 21916
rect 21082 21876 21088 21888
rect 20916 21848 21088 21876
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 21174 21836 21180 21888
rect 21232 21876 21238 21888
rect 23201 21879 23259 21885
rect 23201 21876 23213 21879
rect 21232 21848 23213 21876
rect 21232 21836 21238 21848
rect 23201 21845 23213 21848
rect 23247 21845 23259 21879
rect 23201 21839 23259 21845
rect 23750 21836 23756 21888
rect 23808 21836 23814 21888
rect 24578 21836 24584 21888
rect 24636 21836 24642 21888
rect 24946 21836 24952 21888
rect 25004 21836 25010 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 8846 21672 8852 21684
rect 8619 21644 8852 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 8846 21632 8852 21644
rect 8904 21632 8910 21684
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 9953 21675 10011 21681
rect 9953 21672 9965 21675
rect 9732 21644 9965 21672
rect 9732 21632 9738 21644
rect 9953 21641 9965 21644
rect 9999 21641 10011 21675
rect 9953 21635 10011 21641
rect 10410 21632 10416 21684
rect 10468 21632 10474 21684
rect 10873 21675 10931 21681
rect 10873 21641 10885 21675
rect 10919 21672 10931 21675
rect 10919 21644 12296 21672
rect 10919 21641 10931 21644
rect 10873 21635 10931 21641
rect 8662 21604 8668 21616
rect 6840 21576 8668 21604
rect 4706 21496 4712 21548
rect 4764 21536 4770 21548
rect 6840 21545 6868 21576
rect 8662 21564 8668 21576
rect 8720 21564 8726 21616
rect 11974 21604 11980 21616
rect 9324 21576 11980 21604
rect 5445 21539 5503 21545
rect 5445 21536 5457 21539
rect 4764 21508 5457 21536
rect 4764 21496 4770 21508
rect 5445 21505 5457 21508
rect 5491 21505 5503 21539
rect 5445 21499 5503 21505
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 7466 21496 7472 21548
rect 7524 21536 7530 21548
rect 9324 21545 9352 21576
rect 11974 21564 11980 21576
rect 12032 21564 12038 21616
rect 12268 21604 12296 21644
rect 15102 21632 15108 21684
rect 15160 21672 15166 21684
rect 15749 21675 15807 21681
rect 15160 21644 15516 21672
rect 15160 21632 15166 21644
rect 12802 21604 12808 21616
rect 12268 21576 12808 21604
rect 12802 21564 12808 21576
rect 12860 21564 12866 21616
rect 13170 21564 13176 21616
rect 13228 21564 13234 21616
rect 14458 21604 14464 21616
rect 14398 21576 14464 21604
rect 14458 21564 14464 21576
rect 14516 21604 14522 21616
rect 14642 21604 14648 21616
rect 14516 21576 14648 21604
rect 14516 21564 14522 21576
rect 14642 21564 14648 21576
rect 14700 21564 14706 21616
rect 15488 21604 15516 21644
rect 15749 21641 15761 21675
rect 15795 21672 15807 21675
rect 16666 21672 16672 21684
rect 15795 21644 16672 21672
rect 15795 21641 15807 21644
rect 15749 21635 15807 21641
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 19610 21672 19616 21684
rect 18656 21644 19616 21672
rect 18656 21632 18662 21644
rect 19610 21632 19616 21644
rect 19668 21672 19674 21684
rect 19797 21675 19855 21681
rect 19797 21672 19809 21675
rect 19668 21644 19809 21672
rect 19668 21632 19674 21644
rect 19797 21641 19809 21644
rect 19843 21641 19855 21675
rect 19797 21635 19855 21641
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 21358 21672 21364 21684
rect 20864 21644 21364 21672
rect 20864 21632 20870 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 25409 21675 25467 21681
rect 25409 21672 25421 21675
rect 22388 21644 25421 21672
rect 16025 21607 16083 21613
rect 16025 21604 16037 21607
rect 15488 21576 16037 21604
rect 16025 21573 16037 21576
rect 16071 21604 16083 21607
rect 17126 21604 17132 21616
rect 16071 21576 17132 21604
rect 16071 21573 16083 21576
rect 16025 21567 16083 21573
rect 17126 21564 17132 21576
rect 17184 21564 17190 21616
rect 19153 21607 19211 21613
rect 19153 21573 19165 21607
rect 19199 21604 19211 21607
rect 19702 21604 19708 21616
rect 19199 21576 19708 21604
rect 19199 21573 19211 21576
rect 19153 21567 19211 21573
rect 19702 21564 19708 21576
rect 19760 21564 19766 21616
rect 21082 21564 21088 21616
rect 21140 21604 21146 21616
rect 21450 21604 21456 21616
rect 21140 21576 21456 21604
rect 21140 21564 21146 21576
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 22186 21564 22192 21616
rect 22244 21604 22250 21616
rect 22388 21613 22416 21644
rect 25409 21641 25421 21644
rect 25455 21641 25467 21675
rect 25409 21635 25467 21641
rect 22373 21607 22431 21613
rect 22373 21604 22385 21607
rect 22244 21576 22385 21604
rect 22244 21564 22250 21576
rect 22373 21573 22385 21576
rect 22419 21573 22431 21607
rect 22373 21567 22431 21573
rect 22462 21564 22468 21616
rect 22520 21564 22526 21616
rect 25317 21607 25375 21613
rect 25317 21604 25329 21607
rect 24702 21576 25329 21604
rect 25317 21573 25329 21576
rect 25363 21604 25375 21607
rect 25590 21604 25596 21616
rect 25363 21576 25596 21604
rect 25363 21573 25375 21576
rect 25317 21567 25375 21573
rect 25590 21564 25596 21576
rect 25648 21564 25654 21616
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7524 21508 7941 21536
rect 7524 21496 7530 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 5169 21471 5227 21477
rect 5169 21437 5181 21471
rect 5215 21437 5227 21471
rect 5169 21431 5227 21437
rect 5184 21400 5212 21431
rect 6457 21403 6515 21409
rect 6457 21400 6469 21403
rect 5184 21372 6469 21400
rect 6457 21369 6469 21372
rect 6503 21400 6515 21403
rect 10686 21400 10692 21412
rect 6503 21372 10692 21400
rect 6503 21369 6515 21372
rect 6457 21363 6515 21369
rect 10686 21360 10692 21372
rect 10744 21360 10750 21412
rect 6822 21292 6828 21344
rect 6880 21332 6886 21344
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 6880 21304 7481 21332
rect 6880 21292 6886 21304
rect 7469 21301 7481 21304
rect 7515 21301 7527 21335
rect 10796 21332 10824 21499
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 11112 21508 12081 21536
rect 11112 21496 11118 21508
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21536 15163 21539
rect 16114 21536 16120 21548
rect 15151 21508 16120 21536
rect 15151 21505 15163 21508
rect 15105 21499 15163 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16850 21496 16856 21548
rect 16908 21496 16914 21548
rect 18966 21536 18972 21548
rect 18262 21508 18972 21536
rect 18966 21496 18972 21508
rect 19024 21536 19030 21548
rect 20162 21536 20168 21548
rect 19024 21508 20168 21536
rect 19024 21496 19030 21508
rect 20162 21496 20168 21508
rect 20220 21496 20226 21548
rect 20254 21496 20260 21548
rect 20312 21496 20318 21548
rect 20438 21496 20444 21548
rect 20496 21536 20502 21548
rect 22002 21536 22008 21548
rect 20496 21508 22008 21536
rect 20496 21496 20502 21508
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22278 21536 22284 21548
rect 22152 21508 22284 21536
rect 22152 21496 22158 21508
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 12161 21471 12219 21477
rect 12161 21468 12173 21471
rect 11072 21440 12173 21468
rect 10870 21360 10876 21412
rect 10928 21400 10934 21412
rect 11072 21400 11100 21440
rect 12161 21437 12173 21440
rect 12207 21437 12219 21471
rect 12161 21431 12219 21437
rect 12250 21428 12256 21480
rect 12308 21428 12314 21480
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12406 21440 12909 21468
rect 12406 21412 12434 21440
rect 12897 21437 12909 21440
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 18598 21468 18604 21480
rect 17175 21440 18604 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 20806 21468 20812 21480
rect 19116 21440 20812 21468
rect 19116 21428 19122 21440
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21468 21327 21471
rect 22462 21468 22468 21480
rect 21315 21440 22468 21468
rect 21315 21437 21327 21440
rect 21269 21431 21327 21437
rect 22462 21428 22468 21440
rect 22520 21428 22526 21480
rect 22557 21471 22615 21477
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 22557 21431 22615 21437
rect 10928 21372 11100 21400
rect 10928 21360 10934 21372
rect 11238 21360 11244 21412
rect 11296 21400 11302 21412
rect 12342 21400 12348 21412
rect 11296 21372 12348 21400
rect 11296 21360 11302 21372
rect 12342 21360 12348 21372
rect 12400 21372 12434 21412
rect 18156 21372 22232 21400
rect 12400 21360 12406 21372
rect 11606 21332 11612 21344
rect 10796 21304 11612 21332
rect 7469 21295 7527 21301
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 11701 21335 11759 21341
rect 11701 21301 11713 21335
rect 11747 21332 11759 21335
rect 14182 21332 14188 21344
rect 11747 21304 14188 21332
rect 11747 21301 11759 21304
rect 11701 21295 11759 21301
rect 14182 21292 14188 21304
rect 14240 21292 14246 21344
rect 14642 21292 14648 21344
rect 14700 21292 14706 21344
rect 16298 21292 16304 21344
rect 16356 21292 16362 21344
rect 16390 21292 16396 21344
rect 16448 21332 16454 21344
rect 16485 21335 16543 21341
rect 16485 21332 16497 21335
rect 16448 21304 16497 21332
rect 16448 21292 16454 21304
rect 16485 21301 16497 21304
rect 16531 21332 16543 21335
rect 18156 21332 18184 21372
rect 16531 21304 18184 21332
rect 18601 21335 18659 21341
rect 16531 21301 16543 21304
rect 16485 21295 16543 21301
rect 18601 21301 18613 21335
rect 18647 21332 18659 21335
rect 18782 21332 18788 21344
rect 18647 21304 18788 21332
rect 18647 21301 18659 21304
rect 18601 21295 18659 21301
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 19245 21335 19303 21341
rect 19245 21301 19257 21335
rect 19291 21332 19303 21335
rect 19426 21332 19432 21344
rect 19291 21304 19432 21332
rect 19291 21301 19303 21304
rect 19245 21295 19303 21301
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 20956 21304 22017 21332
rect 20956 21292 20962 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22204 21332 22232 21372
rect 22278 21360 22284 21412
rect 22336 21400 22342 21412
rect 22572 21400 22600 21431
rect 23198 21428 23204 21480
rect 23256 21428 23262 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 24210 21468 24216 21480
rect 23523 21440 24216 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 24210 21428 24216 21440
rect 24268 21428 24274 21480
rect 22336 21372 22600 21400
rect 22336 21360 22342 21372
rect 24026 21332 24032 21344
rect 22204 21304 24032 21332
rect 22005 21295 22063 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24486 21292 24492 21344
rect 24544 21332 24550 21344
rect 24949 21335 25007 21341
rect 24949 21332 24961 21335
rect 24544 21304 24961 21332
rect 24544 21292 24550 21304
rect 24949 21301 24961 21304
rect 24995 21301 25007 21335
rect 24949 21295 25007 21301
rect 25498 21292 25504 21344
rect 25556 21332 25562 21344
rect 25866 21332 25872 21344
rect 25556 21304 25872 21332
rect 25556 21292 25562 21304
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 10318 21088 10324 21140
rect 10376 21128 10382 21140
rect 10413 21131 10471 21137
rect 10413 21128 10425 21131
rect 10376 21100 10425 21128
rect 10376 21088 10382 21100
rect 10413 21097 10425 21100
rect 10459 21097 10471 21131
rect 10413 21091 10471 21097
rect 10686 21088 10692 21140
rect 10744 21128 10750 21140
rect 25130 21128 25136 21140
rect 10744 21100 25136 21128
rect 10744 21088 10750 21100
rect 25130 21088 25136 21100
rect 25188 21128 25194 21140
rect 25498 21128 25504 21140
rect 25188 21100 25504 21128
rect 25188 21088 25194 21100
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 11514 21060 11520 21072
rect 9324 21032 11520 21060
rect 8573 20995 8631 21001
rect 8573 20992 8585 20995
rect 5736 20964 8585 20992
rect 5736 20933 5764 20964
rect 8573 20961 8585 20964
rect 8619 20961 8631 20995
rect 8573 20955 8631 20961
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20893 5779 20927
rect 5721 20887 5779 20893
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 6840 20856 6868 20887
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 7834 20924 7840 20936
rect 7708 20896 7840 20924
rect 7708 20884 7714 20896
rect 7834 20884 7840 20896
rect 7892 20924 7898 20936
rect 9324 20933 9352 21032
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 13354 21020 13360 21072
rect 13412 21060 13418 21072
rect 13538 21060 13544 21072
rect 13412 21032 13544 21060
rect 13412 21020 13418 21032
rect 13538 21020 13544 21032
rect 13596 21020 13602 21072
rect 13909 21063 13967 21069
rect 13909 21029 13921 21063
rect 13955 21060 13967 21063
rect 14918 21060 14924 21072
rect 13955 21032 14924 21060
rect 13955 21029 13967 21032
rect 13909 21023 13967 21029
rect 14918 21020 14924 21032
rect 14976 21020 14982 21072
rect 15286 21020 15292 21072
rect 15344 21020 15350 21072
rect 16390 21020 16396 21072
rect 16448 21020 16454 21072
rect 18598 21020 18604 21072
rect 18656 21020 18662 21072
rect 18966 21020 18972 21072
rect 19024 21020 19030 21072
rect 19429 21063 19487 21069
rect 19429 21029 19441 21063
rect 19475 21060 19487 21063
rect 19702 21060 19708 21072
rect 19475 21032 19708 21060
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 19702 21020 19708 21032
rect 19760 21020 19766 21072
rect 19996 21032 21312 21060
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 10965 20995 11023 21001
rect 10965 20992 10977 20995
rect 9732 20964 10977 20992
rect 9732 20952 9738 20964
rect 10965 20961 10977 20964
rect 11011 20961 11023 20995
rect 10965 20955 11023 20961
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 11609 20995 11667 21001
rect 11609 20992 11621 20995
rect 11296 20964 11621 20992
rect 11296 20952 11302 20964
rect 11609 20961 11621 20964
rect 11655 20961 11667 20995
rect 11609 20955 11667 20961
rect 12618 20952 12624 21004
rect 12676 20992 12682 21004
rect 12676 20964 14688 20992
rect 12676 20952 12682 20964
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7892 20896 7941 20924
rect 7892 20884 7898 20896
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20924 10011 20927
rect 11054 20924 11060 20936
rect 9999 20896 11060 20924
rect 9999 20893 10011 20896
rect 9953 20887 10011 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 14458 20924 14464 20936
rect 13018 20896 14464 20924
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 14660 20933 14688 20964
rect 16298 20952 16304 21004
rect 16356 20992 16362 21004
rect 19996 20992 20024 21032
rect 16356 20964 20024 20992
rect 20073 20995 20131 21001
rect 16356 20952 16362 20964
rect 20073 20961 20085 20995
rect 20119 20992 20131 20995
rect 20346 20992 20352 21004
rect 20119 20964 20352 20992
rect 20119 20961 20131 20964
rect 20073 20955 20131 20961
rect 20346 20952 20352 20964
rect 20404 20952 20410 21004
rect 21284 21001 21312 21032
rect 21818 21020 21824 21072
rect 21876 21020 21882 21072
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 22281 21063 22339 21069
rect 22281 21060 22293 21063
rect 22060 21032 22293 21060
rect 22060 21020 22066 21032
rect 22281 21029 22293 21032
rect 22327 21029 22339 21063
rect 22281 21023 22339 21029
rect 24581 21063 24639 21069
rect 24581 21029 24593 21063
rect 24627 21060 24639 21063
rect 24946 21060 24952 21072
rect 24627 21032 24952 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 24946 21020 24952 21032
rect 25004 21020 25010 21072
rect 21269 20995 21327 21001
rect 21269 20961 21281 20995
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 25038 20992 25044 21004
rect 23891 20964 25044 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 15749 20927 15807 20933
rect 15749 20893 15761 20927
rect 15795 20924 15807 20927
rect 16758 20924 16764 20936
rect 15795 20896 16764 20924
rect 15795 20893 15807 20896
rect 15749 20887 15807 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20924 16911 20927
rect 17034 20924 17040 20936
rect 16899 20896 17040 20924
rect 16899 20893 16911 20896
rect 16853 20887 16911 20893
rect 9122 20856 9128 20868
rect 6840 20828 9128 20856
rect 9122 20816 9128 20828
rect 9180 20816 9186 20868
rect 10781 20859 10839 20865
rect 10781 20825 10793 20859
rect 10827 20856 10839 20859
rect 10827 20828 11652 20856
rect 10827 20825 10839 20828
rect 10781 20819 10839 20825
rect 5074 20748 5080 20800
rect 5132 20748 5138 20800
rect 6365 20791 6423 20797
rect 6365 20757 6377 20791
rect 6411 20788 6423 20791
rect 6638 20788 6644 20800
rect 6411 20760 6644 20788
rect 6411 20757 6423 20760
rect 6365 20751 6423 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 7466 20748 7472 20800
rect 7524 20748 7530 20800
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 10744 20760 10885 20788
rect 10744 20748 10750 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 11624 20788 11652 20828
rect 11882 20816 11888 20868
rect 11940 20816 11946 20868
rect 14550 20856 14556 20868
rect 13280 20828 14556 20856
rect 13280 20788 13308 20828
rect 14550 20816 14556 20828
rect 14608 20816 14614 20868
rect 16298 20816 16304 20868
rect 16356 20856 16362 20868
rect 16868 20856 16896 20887
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 17543 20896 17969 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 19610 20884 19616 20936
rect 19668 20924 19674 20936
rect 19889 20927 19947 20933
rect 19889 20924 19901 20927
rect 19668 20896 19901 20924
rect 19668 20884 19674 20896
rect 19889 20893 19901 20896
rect 19935 20893 19947 20927
rect 21284 20924 21312 20955
rect 25038 20952 25044 20964
rect 25096 20952 25102 21004
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 21284 20896 21496 20924
rect 19889 20887 19947 20893
rect 19058 20856 19064 20868
rect 16356 20828 16896 20856
rect 17236 20828 19064 20856
rect 16356 20816 16362 20828
rect 11624 20760 13308 20788
rect 10873 20751 10931 20757
rect 13354 20748 13360 20800
rect 13412 20748 13418 20800
rect 13630 20748 13636 20800
rect 13688 20748 13694 20800
rect 14182 20748 14188 20800
rect 14240 20748 14246 20800
rect 14369 20791 14427 20797
rect 14369 20757 14381 20791
rect 14415 20788 14427 20791
rect 17236 20788 17264 20828
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 19150 20816 19156 20868
rect 19208 20856 19214 20868
rect 21085 20859 21143 20865
rect 21085 20856 21097 20859
rect 19208 20828 21097 20856
rect 19208 20816 19214 20828
rect 21085 20825 21097 20828
rect 21131 20825 21143 20859
rect 21468 20856 21496 20896
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21876 20896 22017 20924
rect 21876 20884 21882 20896
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20924 22891 20927
rect 23750 20924 23756 20936
rect 22879 20896 23756 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 23750 20884 23756 20896
rect 23808 20884 23814 20936
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 25148 20924 25176 20955
rect 23992 20896 25176 20924
rect 23992 20884 23998 20896
rect 23106 20856 23112 20868
rect 21468 20828 23112 20856
rect 21085 20819 21143 20825
rect 23106 20816 23112 20828
rect 23164 20816 23170 20868
rect 23658 20816 23664 20868
rect 23716 20856 23722 20868
rect 25041 20859 25099 20865
rect 25041 20856 25053 20859
rect 23716 20828 25053 20856
rect 23716 20816 23722 20828
rect 25041 20825 25053 20828
rect 25087 20825 25099 20859
rect 25041 20819 25099 20825
rect 14415 20760 17264 20788
rect 14415 20757 14427 20760
rect 14369 20751 14427 20757
rect 17310 20748 17316 20800
rect 17368 20788 17374 20800
rect 17678 20788 17684 20800
rect 17368 20760 17684 20788
rect 17368 20748 17374 20760
rect 17678 20748 17684 20760
rect 17736 20748 17742 20800
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 18874 20788 18880 20800
rect 18656 20760 18880 20788
rect 18656 20748 18662 20760
rect 18874 20748 18880 20760
rect 18932 20748 18938 20800
rect 19242 20748 19248 20800
rect 19300 20788 19306 20800
rect 19797 20791 19855 20797
rect 19797 20788 19809 20791
rect 19300 20760 19809 20788
rect 19300 20748 19306 20760
rect 19797 20757 19809 20760
rect 19843 20788 19855 20791
rect 20438 20788 20444 20800
rect 19843 20760 20444 20788
rect 19843 20757 19855 20760
rect 19797 20751 19855 20757
rect 20438 20748 20444 20760
rect 20496 20748 20502 20800
rect 20622 20748 20628 20800
rect 20680 20748 20686 20800
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 20993 20791 21051 20797
rect 20993 20788 21005 20791
rect 20864 20760 21005 20788
rect 20864 20748 20870 20760
rect 20993 20757 21005 20760
rect 21039 20757 21051 20791
rect 20993 20751 21051 20757
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 21818 20788 21824 20800
rect 21508 20760 21824 20788
rect 21508 20748 21514 20760
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 24578 20748 24584 20800
rect 24636 20788 24642 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24636 20760 24961 20788
rect 24636 20748 24642 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 5997 20587 6055 20593
rect 5997 20553 6009 20587
rect 6043 20584 6055 20587
rect 6730 20584 6736 20596
rect 6043 20556 6736 20584
rect 6043 20553 6055 20556
rect 5997 20547 6055 20553
rect 6730 20544 6736 20556
rect 6788 20544 6794 20596
rect 10594 20544 10600 20596
rect 10652 20584 10658 20596
rect 10781 20587 10839 20593
rect 10781 20584 10793 20587
rect 10652 20556 10793 20584
rect 10652 20544 10658 20556
rect 10781 20553 10793 20556
rect 10827 20553 10839 20587
rect 10781 20547 10839 20553
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 12345 20587 12403 20593
rect 12345 20584 12357 20587
rect 11940 20556 12357 20584
rect 11940 20544 11946 20556
rect 12345 20553 12357 20556
rect 12391 20553 12403 20587
rect 12345 20547 12403 20553
rect 14642 20544 14648 20596
rect 14700 20544 14706 20596
rect 17586 20544 17592 20596
rect 17644 20584 17650 20596
rect 17644 20556 19104 20584
rect 17644 20544 17650 20556
rect 4893 20519 4951 20525
rect 4893 20485 4905 20519
rect 4939 20516 4951 20519
rect 8110 20516 8116 20528
rect 4939 20488 8116 20516
rect 4939 20485 4951 20488
rect 4893 20479 4951 20485
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 10134 20516 10140 20528
rect 9706 20488 10140 20516
rect 10134 20476 10140 20488
rect 10192 20476 10198 20528
rect 14660 20516 14688 20544
rect 17494 20516 17500 20528
rect 12820 20488 14688 20516
rect 16054 20488 17500 20516
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20448 5411 20451
rect 5994 20448 6000 20460
rect 5399 20420 6000 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 6822 20408 6828 20460
rect 6880 20408 6886 20460
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 8205 20451 8263 20457
rect 8205 20448 8217 20451
rect 7340 20420 8217 20448
rect 7340 20408 7346 20420
rect 8205 20417 8217 20420
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 12820 20457 12848 20488
rect 17494 20476 17500 20488
rect 17552 20516 17558 20528
rect 19076 20516 19104 20556
rect 19150 20544 19156 20596
rect 19208 20544 19214 20596
rect 19334 20544 19340 20596
rect 19392 20544 19398 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 19536 20556 21465 20584
rect 19536 20516 19564 20556
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21600 20556 21833 20584
rect 21600 20544 21606 20556
rect 21821 20553 21833 20556
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 22370 20544 22376 20596
rect 22428 20584 22434 20596
rect 22465 20587 22523 20593
rect 22465 20584 22477 20587
rect 22428 20556 22477 20584
rect 22428 20544 22434 20556
rect 22465 20553 22477 20556
rect 22511 20553 22523 20587
rect 22465 20547 22523 20553
rect 23198 20544 23204 20596
rect 23256 20544 23262 20596
rect 25317 20587 25375 20593
rect 25317 20553 25329 20587
rect 25363 20584 25375 20587
rect 25498 20584 25504 20596
rect 25363 20556 25504 20584
rect 25363 20553 25375 20556
rect 25317 20547 25375 20553
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 22646 20516 22652 20528
rect 17552 20488 17710 20516
rect 19076 20488 19564 20516
rect 20824 20488 22652 20516
rect 17552 20476 17558 20488
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 11112 20420 11713 20448
rect 11112 20408 11118 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 12805 20411 12863 20417
rect 13280 20420 14105 20448
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20380 4399 20383
rect 5074 20380 5080 20392
rect 4387 20352 5080 20380
rect 4387 20349 4399 20352
rect 4341 20343 4399 20349
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 7469 20383 7527 20389
rect 7469 20349 7481 20383
rect 7515 20380 7527 20383
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 7515 20352 8493 20380
rect 7515 20349 7527 20352
rect 7469 20343 7527 20349
rect 8481 20349 8493 20352
rect 8527 20349 8539 20383
rect 8481 20343 8539 20349
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 10229 20383 10287 20389
rect 10229 20380 10241 20383
rect 9180 20352 10241 20380
rect 9180 20340 9186 20352
rect 10229 20349 10241 20352
rect 10275 20380 10287 20383
rect 12250 20380 12256 20392
rect 10275 20352 12256 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 9582 20272 9588 20324
rect 9640 20312 9646 20324
rect 13280 20312 13308 20420
rect 14093 20417 14105 20420
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 16850 20408 16856 20460
rect 16908 20448 16914 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16908 20420 16957 20448
rect 16908 20408 16914 20420
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20714 20448 20720 20460
rect 20027 20420 20720 20448
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 20824 20457 20852 20488
rect 22646 20476 22652 20488
rect 22704 20476 22710 20528
rect 23842 20516 23848 20528
rect 22756 20488 23848 20516
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 21542 20408 21548 20460
rect 21600 20448 21606 20460
rect 22373 20451 22431 20457
rect 22373 20448 22385 20451
rect 21600 20420 22385 20448
rect 21600 20408 21606 20420
rect 22373 20417 22385 20420
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 13722 20340 13728 20392
rect 13780 20380 13786 20392
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 13780 20352 14565 20380
rect 13780 20340 13786 20352
rect 14553 20349 14565 20352
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 14829 20383 14887 20389
rect 14829 20349 14841 20383
rect 14875 20380 14887 20383
rect 16390 20380 16396 20392
rect 14875 20352 16396 20380
rect 14875 20349 14887 20352
rect 14829 20343 14887 20349
rect 16390 20340 16396 20352
rect 16448 20340 16454 20392
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 19242 20380 19248 20392
rect 17267 20352 19248 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 20073 20383 20131 20389
rect 20073 20380 20085 20383
rect 19392 20352 20085 20380
rect 19392 20340 19398 20352
rect 20073 20349 20085 20352
rect 20119 20349 20131 20383
rect 20073 20343 20131 20349
rect 20257 20383 20315 20389
rect 20257 20349 20269 20383
rect 20303 20380 20315 20383
rect 20438 20380 20444 20392
rect 20303 20352 20444 20380
rect 20303 20349 20315 20352
rect 20257 20343 20315 20349
rect 20438 20340 20444 20352
rect 20496 20380 20502 20392
rect 22278 20380 22284 20392
rect 20496 20352 22284 20380
rect 20496 20340 20502 20352
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20380 22707 20383
rect 22756 20380 22784 20488
rect 23842 20476 23848 20488
rect 23900 20476 23906 20528
rect 25130 20516 25136 20528
rect 25070 20488 25136 20516
rect 25130 20476 25136 20488
rect 25188 20476 25194 20528
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23569 20451 23627 20457
rect 23569 20448 23581 20451
rect 23348 20420 23581 20448
rect 23348 20408 23354 20420
rect 23569 20417 23581 20420
rect 23615 20417 23627 20451
rect 23569 20411 23627 20417
rect 22695 20352 22784 20380
rect 22695 20349 22707 20352
rect 22649 20343 22707 20349
rect 9640 20284 13308 20312
rect 9640 20272 9646 20284
rect 22002 20272 22008 20324
rect 22060 20272 22066 20324
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 8570 20244 8576 20256
rect 6972 20216 8576 20244
rect 6972 20204 6978 20216
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 13449 20247 13507 20253
rect 13449 20244 13461 20247
rect 12676 20216 13461 20244
rect 12676 20204 12682 20216
rect 13449 20213 13461 20216
rect 13495 20213 13507 20247
rect 13449 20207 13507 20213
rect 13909 20247 13967 20253
rect 13909 20213 13921 20247
rect 13955 20244 13967 20247
rect 15010 20244 15016 20256
rect 13955 20216 15016 20244
rect 13955 20213 13967 20216
rect 13909 20207 13967 20213
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 15838 20204 15844 20256
rect 15896 20244 15902 20256
rect 16298 20244 16304 20256
rect 15896 20216 16304 20244
rect 15896 20204 15902 20216
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 17678 20204 17684 20256
rect 17736 20244 17742 20256
rect 18693 20247 18751 20253
rect 18693 20244 18705 20247
rect 17736 20216 18705 20244
rect 17736 20204 17742 20216
rect 18693 20213 18705 20216
rect 18739 20213 18751 20247
rect 18693 20207 18751 20213
rect 19610 20204 19616 20256
rect 19668 20204 19674 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 21082 20244 21088 20256
rect 20680 20216 21088 20244
rect 20680 20204 20686 20216
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21542 20204 21548 20256
rect 21600 20244 21606 20256
rect 22664 20244 22692 20343
rect 23842 20340 23848 20392
rect 23900 20340 23906 20392
rect 21600 20216 22692 20244
rect 21600 20204 21606 20216
rect 23106 20204 23112 20256
rect 23164 20244 23170 20256
rect 23658 20244 23664 20256
rect 23164 20216 23664 20244
rect 23164 20204 23170 20216
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7800 20012 7849 20040
rect 7800 20000 7806 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 7837 20003 7895 20009
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 9674 20040 9680 20052
rect 7984 20012 9680 20040
rect 7984 20000 7990 20012
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 9934 20043 9992 20049
rect 9934 20040 9946 20043
rect 9784 20012 9946 20040
rect 6273 19975 6331 19981
rect 6273 19941 6285 19975
rect 6319 19972 6331 19975
rect 9784 19972 9812 20012
rect 9934 20009 9946 20012
rect 9980 20009 9992 20043
rect 9934 20003 9992 20009
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 12894 20040 12900 20052
rect 12584 20012 12900 20040
rect 12584 20000 12590 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13633 20043 13691 20049
rect 13633 20009 13645 20043
rect 13679 20040 13691 20043
rect 16666 20040 16672 20052
rect 13679 20012 16672 20040
rect 13679 20009 13691 20012
rect 13633 20003 13691 20009
rect 6319 19944 9812 19972
rect 6319 19941 6331 19944
rect 6273 19935 6331 19941
rect 12434 19932 12440 19984
rect 12492 19972 12498 19984
rect 12986 19972 12992 19984
rect 12492 19944 12992 19972
rect 12492 19932 12498 19944
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 13648 19972 13676 20003
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16758 20000 16764 20052
rect 16816 20040 16822 20052
rect 17037 20043 17095 20049
rect 17037 20040 17049 20043
rect 16816 20012 17049 20040
rect 16816 20000 16822 20012
rect 17037 20009 17049 20012
rect 17083 20009 17095 20043
rect 17037 20003 17095 20009
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 18230 20040 18236 20052
rect 17552 20012 18236 20040
rect 17552 20000 17558 20012
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 18380 20012 18797 20040
rect 18380 20000 18386 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 18785 20003 18843 20009
rect 13096 19944 13676 19972
rect 18800 19972 18828 20003
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18932 20012 19073 20040
rect 18932 20000 18938 20012
rect 19061 20009 19073 20012
rect 19107 20040 19119 20043
rect 19794 20040 19800 20052
rect 19107 20012 19800 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 22830 20000 22836 20052
rect 22888 20040 22894 20052
rect 25225 20043 25283 20049
rect 25225 20040 25237 20043
rect 22888 20012 25237 20040
rect 22888 20000 22894 20012
rect 25225 20009 25237 20012
rect 25271 20009 25283 20043
rect 25225 20003 25283 20009
rect 18966 19972 18972 19984
rect 18800 19944 18972 19972
rect 4338 19864 4344 19916
rect 4396 19864 4402 19916
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 5644 19876 7389 19904
rect 4614 19796 4620 19848
rect 4672 19796 4678 19848
rect 5644 19845 5672 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 7800 19876 8401 19904
rect 7800 19864 7806 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 9030 19904 9036 19916
rect 8536 19876 9036 19904
rect 8536 19864 8542 19876
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 11146 19904 11152 19916
rect 9692 19876 11152 19904
rect 5629 19839 5687 19845
rect 5629 19805 5641 19839
rect 5675 19805 5687 19839
rect 5629 19799 5687 19805
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6914 19836 6920 19848
rect 6779 19808 6920 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 7282 19796 7288 19848
rect 7340 19836 7346 19848
rect 9692 19845 9720 19876
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 13096 19904 13124 19944
rect 18966 19932 18972 19944
rect 19024 19932 19030 19984
rect 19150 19932 19156 19984
rect 19208 19972 19214 19984
rect 20622 19972 20628 19984
rect 19208 19944 20628 19972
rect 19208 19932 19214 19944
rect 20622 19932 20628 19944
rect 20680 19932 20686 19984
rect 12176 19876 13124 19904
rect 13648 19876 14412 19904
rect 12176 19845 12204 19876
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 7340 19808 9689 19836
rect 7340 19796 7346 19808
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 12161 19839 12219 19845
rect 12161 19805 12173 19839
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 12526 19836 12532 19848
rect 12308 19808 12532 19836
rect 12308 19796 12314 19808
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12618 19796 12624 19848
rect 12676 19796 12682 19848
rect 13648 19836 13676 19876
rect 13556 19808 13676 19836
rect 13909 19839 13967 19845
rect 8205 19771 8263 19777
rect 8205 19737 8217 19771
rect 8251 19768 8263 19771
rect 8251 19740 8432 19768
rect 8251 19737 8263 19740
rect 8205 19731 8263 19737
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 7248 19672 8309 19700
rect 7248 19660 7254 19672
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8404 19700 8432 19740
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 9214 19768 9220 19780
rect 8996 19740 9220 19768
rect 8996 19728 9002 19740
rect 9214 19728 9220 19740
rect 9272 19728 9278 19780
rect 13556 19768 13584 19808
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 13998 19836 14004 19848
rect 13955 19808 14004 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 13998 19796 14004 19808
rect 14056 19836 14062 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14056 19808 14289 19836
rect 14056 19796 14062 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14384 19836 14412 19876
rect 14458 19864 14464 19916
rect 14516 19864 14522 19916
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 14700 19876 15761 19904
rect 14700 19864 14706 19876
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 15749 19867 15807 19873
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 18782 19904 18788 19916
rect 18279 19876 18788 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 18782 19864 18788 19876
rect 18840 19904 18846 19916
rect 18840 19876 19104 19904
rect 18840 19864 18846 19876
rect 15286 19836 15292 19848
rect 14384 19808 15292 19836
rect 14277 19799 14335 19805
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 16393 19839 16451 19845
rect 16393 19805 16405 19839
rect 16439 19836 16451 19839
rect 17494 19836 17500 19848
rect 16439 19808 17500 19836
rect 16439 19805 16451 19808
rect 16393 19799 16451 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19836 18107 19839
rect 18506 19836 18512 19848
rect 18095 19808 18512 19836
rect 18095 19805 18107 19808
rect 18049 19799 18107 19805
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 19076 19836 19104 19876
rect 20070 19864 20076 19916
rect 20128 19904 20134 19916
rect 23845 19907 23903 19913
rect 20128 19876 21864 19904
rect 20128 19864 20134 19876
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 19076 19808 19441 19836
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 20806 19796 20812 19848
rect 20864 19796 20870 19848
rect 10244 19740 10442 19768
rect 11992 19740 13584 19768
rect 8846 19700 8852 19712
rect 8404 19672 8852 19700
rect 8297 19663 8355 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9306 19660 9312 19712
rect 9364 19700 9370 19712
rect 10244 19700 10272 19740
rect 11330 19700 11336 19712
rect 9364 19672 11336 19700
rect 9364 19660 9370 19672
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 11425 19703 11483 19709
rect 11425 19669 11437 19703
rect 11471 19700 11483 19703
rect 11882 19700 11888 19712
rect 11471 19672 11888 19700
rect 11471 19669 11483 19672
rect 11425 19663 11483 19669
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 11992 19709 12020 19740
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 15102 19768 15108 19780
rect 13688 19740 15108 19768
rect 13688 19728 13694 19740
rect 15102 19728 15108 19740
rect 15160 19728 15166 19780
rect 15657 19771 15715 19777
rect 15657 19737 15669 19771
rect 15703 19768 15715 19771
rect 16942 19768 16948 19780
rect 15703 19740 16948 19768
rect 15703 19737 15715 19740
rect 15657 19731 15715 19737
rect 16942 19728 16948 19740
rect 17000 19728 17006 19780
rect 18693 19771 18751 19777
rect 18693 19737 18705 19771
rect 18739 19768 18751 19771
rect 19150 19768 19156 19780
rect 18739 19740 19156 19768
rect 18739 19737 18751 19740
rect 18693 19731 18751 19737
rect 19150 19728 19156 19740
rect 19208 19728 19214 19780
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 21726 19768 21732 19780
rect 19392 19740 21732 19768
rect 19392 19728 19398 19740
rect 21726 19728 21732 19740
rect 21784 19728 21790 19780
rect 11977 19703 12035 19709
rect 11977 19669 11989 19703
rect 12023 19669 12035 19703
rect 11977 19663 12035 19669
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 13265 19703 13323 19709
rect 13265 19700 13277 19703
rect 12308 19672 13277 19700
rect 12308 19660 12314 19672
rect 13265 19669 13277 19672
rect 13311 19669 13323 19703
rect 13265 19663 13323 19669
rect 13906 19660 13912 19712
rect 13964 19700 13970 19712
rect 15197 19703 15255 19709
rect 15197 19700 15209 19703
rect 13964 19672 15209 19700
rect 13964 19660 13970 19672
rect 15197 19669 15209 19672
rect 15243 19669 15255 19703
rect 15197 19663 15255 19669
rect 15562 19660 15568 19712
rect 15620 19660 15626 19712
rect 17586 19660 17592 19712
rect 17644 19660 17650 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18506 19700 18512 19712
rect 18003 19672 18512 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 19058 19660 19064 19712
rect 19116 19700 19122 19712
rect 20073 19703 20131 19709
rect 20073 19700 20085 19703
rect 19116 19672 20085 19700
rect 19116 19660 19122 19672
rect 20073 19669 20085 19672
rect 20119 19669 20131 19703
rect 20073 19663 20131 19669
rect 20346 19660 20352 19712
rect 20404 19660 20410 19712
rect 21836 19700 21864 19876
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24946 19904 24952 19916
rect 23891 19876 24952 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22649 19839 22707 19845
rect 22649 19836 22661 19839
rect 22244 19808 22661 19836
rect 22244 19796 22250 19808
rect 22649 19805 22661 19808
rect 22695 19805 22707 19839
rect 22649 19799 22707 19805
rect 24302 19796 24308 19848
rect 24360 19836 24366 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 24360 19808 24593 19836
rect 24360 19796 24366 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 22005 19771 22063 19777
rect 22005 19737 22017 19771
rect 22051 19768 22063 19771
rect 23382 19768 23388 19780
rect 22051 19740 23388 19768
rect 22051 19737 22063 19740
rect 22005 19731 22063 19737
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 22370 19700 22376 19712
rect 21836 19672 22376 19700
rect 22370 19660 22376 19672
rect 22428 19700 22434 19712
rect 25130 19700 25136 19712
rect 22428 19672 25136 19700
rect 22428 19660 22434 19672
rect 25130 19660 25136 19672
rect 25188 19660 25194 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 4338 19456 4344 19508
rect 4396 19496 4402 19508
rect 4985 19499 5043 19505
rect 4985 19496 4997 19499
rect 4396 19468 4997 19496
rect 4396 19456 4402 19468
rect 4985 19465 4997 19468
rect 5031 19465 5043 19499
rect 4985 19459 5043 19465
rect 5994 19456 6000 19508
rect 6052 19456 6058 19508
rect 6641 19499 6699 19505
rect 6641 19465 6653 19499
rect 6687 19496 6699 19499
rect 8478 19496 8484 19508
rect 6687 19468 8484 19496
rect 6687 19465 6699 19468
rect 6641 19459 6699 19465
rect 8478 19456 8484 19468
rect 8536 19456 8542 19508
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 9033 19499 9091 19505
rect 9033 19496 9045 19499
rect 8628 19468 9045 19496
rect 8628 19456 8634 19468
rect 9033 19465 9045 19468
rect 9079 19465 9091 19499
rect 9033 19459 9091 19465
rect 7834 19428 7840 19440
rect 5368 19400 7840 19428
rect 3970 19320 3976 19372
rect 4028 19320 4034 19372
rect 5368 19369 5396 19400
rect 7834 19388 7840 19400
rect 7892 19388 7898 19440
rect 8294 19388 8300 19440
rect 8352 19388 8358 19440
rect 9048 19428 9076 19459
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 9585 19499 9643 19505
rect 9585 19496 9597 19499
rect 9548 19468 9597 19496
rect 9548 19456 9554 19468
rect 9585 19465 9597 19468
rect 9631 19465 9643 19499
rect 9585 19459 9643 19465
rect 9692 19468 10167 19496
rect 9692 19428 9720 19468
rect 9048 19400 9720 19428
rect 9766 19388 9772 19440
rect 9824 19428 9830 19440
rect 10045 19431 10103 19437
rect 10045 19428 10057 19431
rect 9824 19400 10057 19428
rect 9824 19388 9830 19400
rect 10045 19397 10057 19400
rect 10091 19397 10103 19431
rect 10139 19428 10167 19468
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10468 19468 10977 19496
rect 10468 19456 10474 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 12253 19499 12311 19505
rect 12253 19465 12265 19499
rect 12299 19496 12311 19499
rect 15194 19496 15200 19508
rect 12299 19468 15200 19496
rect 12299 19465 12311 19468
rect 12253 19459 12311 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19465 15899 19499
rect 15841 19459 15899 19465
rect 12066 19428 12072 19440
rect 10139 19400 12072 19428
rect 10045 19391 10103 19397
rect 12066 19388 12072 19400
rect 12124 19388 12130 19440
rect 12986 19428 12992 19440
rect 12636 19400 12992 19428
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 7282 19320 7288 19372
rect 7340 19320 7346 19372
rect 9953 19363 10011 19369
rect 9953 19360 9965 19363
rect 8772 19332 9965 19360
rect 3694 19252 3700 19304
rect 3752 19252 3758 19304
rect 4246 19252 4252 19304
rect 4304 19292 4310 19304
rect 4801 19295 4859 19301
rect 4801 19292 4813 19295
rect 4304 19264 4813 19292
rect 4304 19252 4310 19264
rect 4801 19261 4813 19264
rect 4847 19261 4859 19295
rect 7561 19295 7619 19301
rect 7561 19292 7573 19295
rect 4801 19255 4859 19261
rect 6748 19264 7573 19292
rect 5994 19184 6000 19236
rect 6052 19224 6058 19236
rect 6748 19224 6776 19264
rect 7561 19261 7573 19264
rect 7607 19261 7619 19295
rect 7561 19255 7619 19261
rect 7926 19252 7932 19304
rect 7984 19292 7990 19304
rect 8772 19292 8800 19332
rect 9953 19329 9965 19332
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11422 19360 11428 19372
rect 11195 19332 11428 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12636 19369 12664 19400
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 13538 19388 13544 19440
rect 13596 19428 13602 19440
rect 13596 19400 14858 19428
rect 13596 19388 13602 19400
rect 12621 19363 12679 19369
rect 11940 19332 12434 19360
rect 11940 19320 11946 19332
rect 7984 19264 8800 19292
rect 10229 19295 10287 19301
rect 7984 19252 7990 19264
rect 10229 19261 10241 19295
rect 10275 19292 10287 19295
rect 12406 19292 12434 19332
rect 12621 19329 12633 19363
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 12894 19360 12900 19372
rect 12759 19332 12900 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 13780 19332 14105 19360
rect 13780 19320 13786 19332
rect 14093 19329 14105 19332
rect 14139 19329 14151 19363
rect 15856 19360 15884 19459
rect 17494 19456 17500 19508
rect 17552 19456 17558 19508
rect 17957 19499 18015 19505
rect 17957 19465 17969 19499
rect 18003 19496 18015 19499
rect 19334 19496 19340 19508
rect 18003 19468 19340 19496
rect 18003 19465 18015 19468
rect 17957 19459 18015 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 20622 19496 20628 19508
rect 19720 19468 20628 19496
rect 16206 19388 16212 19440
rect 16264 19428 16270 19440
rect 16264 19400 19288 19428
rect 16264 19388 16270 19400
rect 16390 19360 16396 19372
rect 15856 19332 16396 19360
rect 14093 19323 14151 19329
rect 16390 19320 16396 19332
rect 16448 19360 16454 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16448 19332 16865 19360
rect 16448 19320 16454 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 18141 19363 18199 19369
rect 18141 19329 18153 19363
rect 18187 19360 18199 19363
rect 18414 19360 18420 19372
rect 18187 19332 18420 19360
rect 18187 19329 18199 19332
rect 18141 19323 18199 19329
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19360 18659 19363
rect 19058 19360 19064 19372
rect 18647 19332 19064 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 19260 19360 19288 19400
rect 19334 19360 19340 19372
rect 19260 19332 19340 19360
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19720 19369 19748 19468
rect 20622 19456 20628 19468
rect 20680 19496 20686 19508
rect 22278 19496 22284 19508
rect 20680 19468 22284 19496
rect 20680 19456 20686 19468
rect 20070 19388 20076 19440
rect 20128 19428 20134 19440
rect 22066 19428 22094 19468
rect 22278 19456 22284 19468
rect 22336 19496 22342 19508
rect 23290 19496 23296 19508
rect 22336 19468 23296 19496
rect 22336 19456 22342 19468
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 23750 19456 23756 19508
rect 23808 19496 23814 19508
rect 24213 19499 24271 19505
rect 24213 19496 24225 19499
rect 23808 19468 24225 19496
rect 23808 19456 23814 19468
rect 24213 19465 24225 19468
rect 24259 19465 24271 19499
rect 24213 19459 24271 19465
rect 24670 19456 24676 19508
rect 24728 19456 24734 19508
rect 25498 19456 25504 19508
rect 25556 19456 25562 19508
rect 20128 19400 20470 19428
rect 22020 19400 22094 19428
rect 20128 19388 20134 19400
rect 22020 19369 22048 19400
rect 22370 19388 22376 19440
rect 22428 19428 22434 19440
rect 22428 19400 22770 19428
rect 22428 19388 22434 19400
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19329 22063 19363
rect 23934 19360 23940 19372
rect 22005 19323 22063 19329
rect 23768 19332 23940 19360
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 10275 19264 12112 19292
rect 12406 19264 12817 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 6052 19196 6776 19224
rect 6052 19184 6058 19196
rect 8570 19184 8576 19236
rect 8628 19224 8634 19236
rect 9306 19224 9312 19236
rect 8628 19196 9312 19224
rect 8628 19184 8634 19196
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 2774 19116 2780 19168
rect 2832 19156 2838 19168
rect 8202 19156 8208 19168
rect 2832 19128 8208 19156
rect 2832 19116 2838 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 10594 19116 10600 19168
rect 10652 19116 10658 19168
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 10928 19128 11529 19156
rect 10928 19116 10934 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 11790 19116 11796 19168
rect 11848 19116 11854 19168
rect 11974 19116 11980 19168
rect 12032 19116 12038 19168
rect 12084 19156 12112 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13446 19252 13452 19304
rect 13504 19252 13510 19304
rect 12342 19184 12348 19236
rect 12400 19224 12406 19236
rect 12710 19224 12716 19236
rect 12400 19196 12716 19224
rect 12400 19184 12406 19196
rect 12710 19184 12716 19196
rect 12768 19224 12774 19236
rect 13740 19224 13768 19320
rect 14366 19252 14372 19304
rect 14424 19252 14430 19304
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 18322 19292 18328 19304
rect 15160 19264 18328 19292
rect 15160 19252 15166 19264
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19024 19264 19993 19292
rect 19024 19252 19030 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 22281 19295 22339 19301
rect 22281 19261 22293 19295
rect 22327 19292 22339 19295
rect 22738 19292 22744 19304
rect 22327 19264 22744 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 23768 19301 23796 19332
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 24044 19332 24593 19360
rect 23753 19295 23811 19301
rect 23753 19261 23765 19295
rect 23799 19261 23811 19295
rect 23753 19255 23811 19261
rect 12768 19196 13768 19224
rect 12768 19184 12774 19196
rect 15746 19184 15752 19236
rect 15804 19224 15810 19236
rect 18138 19224 18144 19236
rect 15804 19196 18144 19224
rect 15804 19184 15810 19196
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 18288 19196 19748 19224
rect 18288 19184 18294 19196
rect 14182 19156 14188 19168
rect 12084 19128 14188 19156
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 16206 19156 16212 19168
rect 15436 19128 16212 19156
rect 15436 19116 15442 19128
rect 16206 19116 16212 19128
rect 16264 19116 16270 19168
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 16393 19159 16451 19165
rect 16393 19156 16405 19159
rect 16356 19128 16405 19156
rect 16356 19116 16362 19128
rect 16393 19125 16405 19128
rect 16439 19125 16451 19159
rect 16393 19119 16451 19125
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19245 19159 19303 19165
rect 19245 19156 19257 19159
rect 19116 19128 19257 19156
rect 19116 19116 19122 19128
rect 19245 19125 19257 19128
rect 19291 19125 19303 19159
rect 19720 19156 19748 19196
rect 23474 19184 23480 19236
rect 23532 19224 23538 19236
rect 24044 19233 24072 19332
rect 24581 19329 24593 19332
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 24486 19252 24492 19304
rect 24544 19292 24550 19304
rect 24765 19295 24823 19301
rect 24765 19292 24777 19295
rect 24544 19264 24777 19292
rect 24544 19252 24550 19264
rect 24765 19261 24777 19264
rect 24811 19261 24823 19295
rect 24765 19255 24823 19261
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 25225 19295 25283 19301
rect 25225 19292 25237 19295
rect 25188 19264 25237 19292
rect 25188 19252 25194 19264
rect 25225 19261 25237 19264
rect 25271 19292 25283 19295
rect 26142 19292 26148 19304
rect 25271 19264 26148 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 24029 19227 24087 19233
rect 24029 19224 24041 19227
rect 23532 19196 24041 19224
rect 23532 19184 23538 19196
rect 24029 19193 24041 19196
rect 24075 19193 24087 19227
rect 24029 19187 24087 19193
rect 20070 19156 20076 19168
rect 19720 19128 20076 19156
rect 19245 19119 19303 19125
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 20588 19128 21465 19156
rect 20588 19116 20594 19128
rect 21453 19125 21465 19128
rect 21499 19125 21511 19159
rect 21453 19119 21511 19125
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 13906 18952 13912 18964
rect 4908 18924 13912 18952
rect 4246 18708 4252 18760
rect 4304 18708 4310 18760
rect 4908 18757 4936 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 15010 18912 15016 18964
rect 15068 18952 15074 18964
rect 15068 18924 20208 18952
rect 15068 18912 15074 18924
rect 5994 18844 6000 18896
rect 6052 18844 6058 18896
rect 9582 18844 9588 18896
rect 9640 18844 9646 18896
rect 10781 18887 10839 18893
rect 10781 18853 10793 18887
rect 10827 18884 10839 18887
rect 11330 18884 11336 18896
rect 10827 18856 11336 18884
rect 10827 18853 10839 18856
rect 10781 18847 10839 18853
rect 11330 18844 11336 18856
rect 11388 18844 11394 18896
rect 16390 18844 16396 18896
rect 16448 18884 16454 18896
rect 16448 18856 16620 18884
rect 16448 18844 16454 18856
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7282 18816 7288 18828
rect 6687 18788 7288 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 8110 18816 8116 18828
rect 8036 18788 8116 18816
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18717 4951 18751
rect 4893 18711 4951 18717
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5994 18748 6000 18760
rect 5399 18720 6000 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 8036 18748 8064 18788
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 8444 18788 10149 18816
rect 8444 18776 8450 18788
rect 10137 18785 10149 18788
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 10594 18776 10600 18828
rect 10652 18816 10658 18828
rect 11241 18819 11299 18825
rect 11241 18816 11253 18819
rect 10652 18788 11253 18816
rect 10652 18776 10658 18788
rect 11241 18785 11253 18788
rect 11287 18785 11299 18819
rect 11241 18779 11299 18785
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18816 11483 18819
rect 11698 18816 11704 18828
rect 11471 18788 11704 18816
rect 11471 18785 11483 18788
rect 11425 18779 11483 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12342 18816 12348 18828
rect 12023 18788 12348 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 14458 18776 14464 18828
rect 14516 18816 14522 18828
rect 14516 18788 16436 18816
rect 14516 18776 14522 18788
rect 8570 18748 8576 18760
rect 8036 18734 8576 18748
rect 8050 18720 8576 18734
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9953 18751 10011 18757
rect 9953 18748 9965 18751
rect 8720 18720 9965 18748
rect 8720 18708 8726 18720
rect 9953 18717 9965 18720
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 11054 18748 11060 18760
rect 10091 18720 11060 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13740 18720 14289 18748
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 3237 18683 3295 18689
rect 3237 18680 3249 18683
rect 3191 18652 3249 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3237 18649 3249 18652
rect 3283 18680 3295 18683
rect 3283 18652 6224 18680
rect 3283 18649 3295 18652
rect 3237 18643 3295 18649
rect 4062 18572 4068 18624
rect 4120 18572 4126 18624
rect 4522 18572 4528 18624
rect 4580 18612 4586 18624
rect 4709 18615 4767 18621
rect 4709 18612 4721 18615
rect 4580 18584 4721 18612
rect 4580 18572 4586 18584
rect 4709 18581 4721 18584
rect 4755 18581 4767 18615
rect 6196 18612 6224 18652
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 6917 18683 6975 18689
rect 6917 18680 6929 18683
rect 6696 18652 6929 18680
rect 6696 18640 6702 18652
rect 6917 18649 6929 18652
rect 6963 18649 6975 18683
rect 12158 18680 12164 18692
rect 6917 18643 6975 18649
rect 8220 18652 12164 18680
rect 8220 18612 8248 18652
rect 12158 18640 12164 18652
rect 12216 18640 12222 18692
rect 12250 18640 12256 18692
rect 12308 18640 12314 18692
rect 13538 18680 13544 18692
rect 13478 18652 13544 18680
rect 13538 18640 13544 18652
rect 13596 18640 13602 18692
rect 6196 18584 8248 18612
rect 4709 18575 4767 18581
rect 9030 18572 9036 18624
rect 9088 18572 9094 18624
rect 9214 18572 9220 18624
rect 9272 18572 9278 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11149 18615 11207 18621
rect 11149 18612 11161 18615
rect 11112 18584 11161 18612
rect 11112 18572 11118 18584
rect 11149 18581 11161 18584
rect 11195 18581 11207 18615
rect 11149 18575 11207 18581
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 12066 18612 12072 18624
rect 11388 18584 12072 18612
rect 11388 18572 11394 18584
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 13556 18612 13584 18640
rect 12400 18584 13584 18612
rect 12400 18572 12406 18584
rect 13630 18572 13636 18624
rect 13688 18612 13694 18624
rect 13740 18621 13768 18720
rect 14277 18717 14289 18720
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 16408 18757 16436 18788
rect 16482 18776 16488 18828
rect 16540 18776 16546 18828
rect 16592 18825 16620 18856
rect 18138 18844 18144 18896
rect 18196 18844 18202 18896
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 18782 18884 18788 18896
rect 18380 18856 18788 18884
rect 18380 18844 18386 18856
rect 18782 18844 18788 18856
rect 18840 18884 18846 18896
rect 18877 18887 18935 18893
rect 18877 18884 18889 18887
rect 18840 18856 18889 18884
rect 18840 18844 18846 18856
rect 18877 18853 18889 18856
rect 18923 18853 18935 18887
rect 18877 18847 18935 18853
rect 16577 18819 16635 18825
rect 16577 18785 16589 18819
rect 16623 18785 16635 18819
rect 20180 18816 20208 18924
rect 20254 18912 20260 18964
rect 20312 18952 20318 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 20312 18924 21465 18952
rect 20312 18912 20318 18924
rect 21453 18921 21465 18924
rect 21499 18921 21511 18955
rect 21453 18915 21511 18921
rect 21910 18912 21916 18964
rect 21968 18912 21974 18964
rect 25225 18955 25283 18961
rect 25225 18921 25237 18955
rect 25271 18952 25283 18955
rect 26050 18952 26056 18964
rect 25271 18924 26056 18952
rect 25271 18921 25283 18924
rect 25225 18915 25283 18921
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 20530 18844 20536 18896
rect 20588 18884 20594 18896
rect 20588 18856 20852 18884
rect 20588 18844 20594 18856
rect 20824 18825 20852 18856
rect 20809 18819 20867 18825
rect 20180 18788 20760 18816
rect 16577 18779 16635 18785
rect 15565 18751 15623 18757
rect 15565 18748 15577 18751
rect 15252 18720 15577 18748
rect 15252 18708 15258 18720
rect 15565 18717 15577 18720
rect 15611 18717 15623 18751
rect 15565 18711 15623 18717
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17770 18748 17776 18760
rect 17267 18720 17776 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 17880 18720 19533 18748
rect 17880 18680 17908 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 19668 18720 20545 18748
rect 19668 18708 19674 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20732 18748 20760 18788
rect 20809 18785 20821 18819
rect 20855 18785 20867 18819
rect 20809 18779 20867 18785
rect 22278 18776 22284 18828
rect 22336 18776 22342 18828
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 23624 18788 24624 18816
rect 23624 18776 23630 18788
rect 24596 18757 24624 18788
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 20732 18720 21649 18748
rect 20533 18711 20591 18717
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 15396 18652 17908 18680
rect 18693 18683 18751 18689
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13688 18584 13737 18612
rect 13688 18572 13694 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 13725 18575 13783 18581
rect 14921 18615 14979 18621
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15010 18612 15016 18624
rect 14967 18584 15016 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15396 18621 15424 18652
rect 18693 18649 18705 18683
rect 18739 18680 18751 18683
rect 18874 18680 18880 18692
rect 18739 18652 18880 18680
rect 18739 18649 18751 18652
rect 18693 18643 18751 18649
rect 18874 18640 18880 18652
rect 18932 18640 18938 18692
rect 19705 18683 19763 18689
rect 19705 18649 19717 18683
rect 19751 18680 19763 18683
rect 22186 18680 22192 18692
rect 19751 18652 22192 18680
rect 19751 18649 19763 18652
rect 19705 18643 19763 18649
rect 22186 18640 22192 18652
rect 22244 18640 22250 18692
rect 22278 18640 22284 18692
rect 22336 18680 22342 18692
rect 22557 18683 22615 18689
rect 22557 18680 22569 18683
rect 22336 18652 22569 18680
rect 22336 18640 22342 18652
rect 22557 18649 22569 18652
rect 22603 18649 22615 18683
rect 22557 18643 22615 18649
rect 22664 18652 23046 18680
rect 15381 18615 15439 18621
rect 15381 18581 15393 18615
rect 15427 18581 15439 18615
rect 15381 18575 15439 18581
rect 16022 18572 16028 18624
rect 16080 18572 16086 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17865 18615 17923 18621
rect 17865 18612 17877 18615
rect 17184 18584 17877 18612
rect 17184 18572 17190 18584
rect 17865 18581 17877 18584
rect 17911 18581 17923 18615
rect 17865 18575 17923 18581
rect 20162 18572 20168 18624
rect 20220 18572 20226 18624
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18612 20683 18615
rect 20898 18612 20904 18624
rect 20671 18584 20904 18612
rect 20671 18581 20683 18584
rect 20625 18575 20683 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 22370 18572 22376 18624
rect 22428 18612 22434 18624
rect 22664 18612 22692 18652
rect 22428 18584 22692 18612
rect 22428 18572 22434 18584
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 24029 18615 24087 18621
rect 24029 18612 24041 18615
rect 23624 18584 24041 18612
rect 23624 18572 23630 18584
rect 24029 18581 24041 18584
rect 24075 18581 24087 18615
rect 24029 18575 24087 18581
rect 24210 18572 24216 18624
rect 24268 18612 24274 18624
rect 25498 18612 25504 18624
rect 24268 18584 25504 18612
rect 24268 18572 24274 18584
rect 25498 18572 25504 18584
rect 25556 18572 25562 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 5994 18368 6000 18420
rect 6052 18368 6058 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 9769 18411 9827 18417
rect 9769 18408 9781 18411
rect 9732 18380 9781 18408
rect 9732 18368 9738 18380
rect 9769 18377 9781 18380
rect 9815 18408 9827 18411
rect 10318 18408 10324 18420
rect 9815 18380 10324 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 10502 18408 10508 18420
rect 10459 18380 10508 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 12345 18411 12403 18417
rect 12345 18408 12357 18411
rect 11572 18380 12357 18408
rect 11572 18368 11578 18380
rect 12345 18377 12357 18380
rect 12391 18377 12403 18411
rect 12345 18371 12403 18377
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18377 12955 18411
rect 12897 18371 12955 18377
rect 13265 18411 13323 18417
rect 13265 18377 13277 18411
rect 13311 18408 13323 18411
rect 13446 18408 13452 18420
rect 13311 18380 13452 18408
rect 13311 18377 13323 18380
rect 13265 18371 13323 18377
rect 4522 18300 4528 18352
rect 4580 18300 4586 18352
rect 8386 18340 8392 18352
rect 6932 18312 8392 18340
rect 6932 18281 6960 18312
rect 8386 18300 8392 18312
rect 8444 18300 8450 18352
rect 8570 18300 8576 18352
rect 8628 18340 8634 18352
rect 8628 18312 8786 18340
rect 8628 18300 8634 18312
rect 9950 18300 9956 18352
rect 10008 18340 10014 18352
rect 10045 18343 10103 18349
rect 10045 18340 10057 18343
rect 10008 18312 10057 18340
rect 10008 18300 10014 18312
rect 10045 18309 10057 18312
rect 10091 18340 10103 18343
rect 10781 18343 10839 18349
rect 10781 18340 10793 18343
rect 10091 18312 10793 18340
rect 10091 18309 10103 18312
rect 10045 18303 10103 18309
rect 10781 18309 10793 18312
rect 10827 18309 10839 18343
rect 10781 18303 10839 18309
rect 10873 18343 10931 18349
rect 10873 18309 10885 18343
rect 10919 18340 10931 18343
rect 12802 18340 12808 18352
rect 10919 18312 12808 18340
rect 10919 18309 10931 18312
rect 10873 18303 10931 18309
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 12912 18340 12940 18371
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14424 18380 15209 18408
rect 14424 18368 14430 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 19242 18368 19248 18420
rect 19300 18408 19306 18420
rect 19705 18411 19763 18417
rect 19705 18408 19717 18411
rect 19300 18380 19717 18408
rect 19300 18368 19306 18380
rect 19705 18377 19717 18380
rect 19751 18377 19763 18411
rect 19705 18371 19763 18377
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20165 18411 20223 18417
rect 20165 18408 20177 18411
rect 20036 18380 20177 18408
rect 20036 18368 20042 18380
rect 20165 18377 20177 18380
rect 20211 18377 20223 18411
rect 20165 18371 20223 18377
rect 21453 18411 21511 18417
rect 21453 18377 21465 18411
rect 21499 18408 21511 18411
rect 22094 18408 22100 18420
rect 21499 18380 22100 18408
rect 21499 18377 21511 18380
rect 21453 18371 21511 18377
rect 22094 18368 22100 18380
rect 22152 18368 22158 18420
rect 13814 18340 13820 18352
rect 12912 18312 13820 18340
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 14826 18300 14832 18352
rect 14884 18340 14890 18352
rect 16301 18343 16359 18349
rect 16301 18340 16313 18343
rect 14884 18312 16313 18340
rect 14884 18300 14890 18312
rect 16301 18309 16313 18312
rect 16347 18309 16359 18343
rect 16301 18303 16359 18309
rect 17126 18300 17132 18352
rect 17184 18300 17190 18352
rect 18414 18340 18420 18352
rect 18354 18312 18420 18340
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 18598 18300 18604 18352
rect 18656 18340 18662 18352
rect 18656 18312 22048 18340
rect 18656 18300 18662 18312
rect 3973 18275 4031 18281
rect 3973 18241 3985 18275
rect 4019 18241 4031 18275
rect 3973 18235 4031 18241
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18241 5411 18275
rect 5353 18235 5411 18241
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 3786 18028 3792 18080
rect 3844 18028 3850 18080
rect 3988 18068 4016 18235
rect 4706 18164 4712 18216
rect 4764 18164 4770 18216
rect 5368 18204 5396 18235
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7340 18244 8033 18272
rect 7340 18232 7346 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 11422 18272 11428 18284
rect 8021 18235 8079 18241
rect 10980 18244 11428 18272
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 5368 18176 7573 18204
rect 7561 18173 7573 18176
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18204 8355 18207
rect 10980 18204 11008 18244
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 11882 18272 11888 18284
rect 11747 18244 11888 18272
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 14553 18275 14611 18281
rect 12216 18244 14504 18272
rect 12216 18232 12222 18244
rect 8343 18176 11008 18204
rect 11057 18207 11115 18213
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 11057 18173 11069 18207
rect 11103 18204 11115 18207
rect 12066 18204 12072 18216
rect 11103 18176 12072 18204
rect 11103 18173 11115 18176
rect 11057 18167 11115 18173
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 13354 18164 13360 18216
rect 13412 18164 13418 18216
rect 13446 18164 13452 18216
rect 13504 18164 13510 18216
rect 14476 18204 14504 18244
rect 14553 18241 14565 18275
rect 14599 18272 14611 18275
rect 15286 18272 15292 18284
rect 14599 18244 15292 18272
rect 14599 18241 14611 18244
rect 14553 18235 14611 18241
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15528 18244 15669 18272
rect 15528 18232 15534 18244
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 18432 18272 18460 18300
rect 18874 18272 18880 18284
rect 18432 18244 18880 18272
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 19058 18232 19064 18284
rect 19116 18232 19122 18284
rect 22020 18281 22048 18312
rect 22370 18300 22376 18352
rect 22428 18340 22434 18352
rect 22428 18312 24242 18340
rect 22428 18300 22434 18312
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 20824 18204 20852 18235
rect 23290 18232 23296 18284
rect 23348 18272 23354 18284
rect 23477 18275 23535 18281
rect 23477 18272 23489 18275
rect 23348 18244 23489 18272
rect 23348 18232 23354 18244
rect 23477 18241 23489 18244
rect 23523 18241 23535 18275
rect 23477 18235 23535 18241
rect 22649 18207 22707 18213
rect 22649 18204 22661 18207
rect 14476 18176 19196 18204
rect 20824 18176 22661 18204
rect 16022 18136 16028 18148
rect 9324 18108 16028 18136
rect 9324 18068 9352 18108
rect 16022 18096 16028 18108
rect 16080 18096 16086 18148
rect 19168 18136 19196 18176
rect 22649 18173 22661 18176
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 23753 18207 23811 18213
rect 23753 18173 23765 18207
rect 23799 18204 23811 18207
rect 25590 18204 25596 18216
rect 23799 18176 25596 18204
rect 23799 18173 23811 18176
rect 23753 18167 23811 18173
rect 25590 18164 25596 18176
rect 25648 18164 25654 18216
rect 22002 18136 22008 18148
rect 19168 18108 22008 18136
rect 22002 18096 22008 18108
rect 22060 18136 22066 18148
rect 23474 18136 23480 18148
rect 22060 18108 23480 18136
rect 22060 18096 22066 18108
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 3988 18040 9352 18068
rect 13906 18028 13912 18080
rect 13964 18028 13970 18080
rect 14182 18028 14188 18080
rect 14240 18028 14246 18080
rect 18598 18028 18604 18080
rect 18656 18028 18662 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 22094 18068 22100 18080
rect 20220 18040 22100 18068
rect 20220 18028 20226 18040
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 22830 18028 22836 18080
rect 22888 18068 22894 18080
rect 23017 18071 23075 18077
rect 23017 18068 23029 18071
rect 22888 18040 23029 18068
rect 22888 18028 22894 18040
rect 23017 18037 23029 18040
rect 23063 18037 23075 18071
rect 23017 18031 23075 18037
rect 25130 18028 25136 18080
rect 25188 18068 25194 18080
rect 25225 18071 25283 18077
rect 25225 18068 25237 18071
rect 25188 18040 25237 18068
rect 25188 18028 25194 18040
rect 25225 18037 25237 18040
rect 25271 18037 25283 18071
rect 25225 18031 25283 18037
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 7834 17864 7840 17876
rect 3252 17836 7840 17864
rect 3252 17737 3280 17836
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 9125 17867 9183 17873
rect 9125 17833 9137 17867
rect 9171 17864 9183 17867
rect 9306 17864 9312 17876
rect 9171 17836 9312 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 10962 17864 10968 17876
rect 9416 17836 10968 17864
rect 5169 17799 5227 17805
rect 5169 17765 5181 17799
rect 5215 17796 5227 17799
rect 9416 17796 9444 17836
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 11330 17824 11336 17876
rect 11388 17864 11394 17876
rect 12158 17864 12164 17876
rect 11388 17836 12164 17864
rect 11388 17824 11394 17836
rect 12158 17824 12164 17836
rect 12216 17864 12222 17876
rect 12342 17864 12348 17876
rect 12216 17836 12348 17864
rect 12216 17824 12222 17836
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12860 17836 13001 17864
rect 12860 17824 12866 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 13262 17824 13268 17876
rect 13320 17864 13326 17876
rect 15194 17864 15200 17876
rect 13320 17836 15200 17864
rect 13320 17824 13326 17836
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 15286 17824 15292 17876
rect 15344 17824 15350 17876
rect 15746 17824 15752 17876
rect 15804 17824 15810 17876
rect 20990 17824 20996 17876
rect 21048 17864 21054 17876
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 21048 17836 21097 17864
rect 21048 17824 21054 17836
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 22189 17867 22247 17873
rect 22189 17864 22201 17867
rect 21085 17827 21143 17833
rect 21192 17836 22201 17864
rect 5215 17768 5764 17796
rect 5215 17765 5227 17768
rect 5169 17759 5227 17765
rect 3237 17731 3295 17737
rect 3237 17697 3249 17731
rect 3283 17697 3295 17731
rect 3237 17691 3295 17697
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 5442 17728 5448 17740
rect 4295 17700 5448 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 4724 17669 4752 17700
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17660 5411 17663
rect 5626 17660 5632 17672
rect 5399 17632 5632 17660
rect 5399 17629 5411 17632
rect 5353 17623 5411 17629
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 5736 17660 5764 17768
rect 5828 17768 9444 17796
rect 5828 17737 5856 17768
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 12492 17768 13584 17796
rect 12492 17756 12498 17768
rect 5813 17731 5871 17737
rect 5813 17697 5825 17731
rect 5859 17697 5871 17731
rect 5813 17691 5871 17697
rect 6454 17688 6460 17740
rect 6512 17688 6518 17740
rect 7742 17728 7748 17740
rect 6840 17700 7748 17728
rect 6840 17669 6868 17700
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9180 17700 9689 17728
rect 9180 17688 9186 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 10781 17731 10839 17737
rect 10781 17728 10793 17731
rect 9677 17691 9735 17697
rect 9784 17700 10793 17728
rect 6825 17663 6883 17669
rect 5736 17632 6776 17660
rect 6365 17595 6423 17601
rect 6365 17561 6377 17595
rect 6411 17592 6423 17595
rect 6546 17592 6552 17604
rect 6411 17564 6552 17592
rect 6411 17561 6423 17564
rect 6365 17555 6423 17561
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 6748 17592 6776 17632
rect 6825 17629 6837 17663
rect 6871 17629 6883 17663
rect 6825 17623 6883 17629
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7524 17632 7941 17660
rect 7524 17620 7530 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 9784 17660 9812 17700
rect 10781 17697 10793 17700
rect 10827 17697 10839 17731
rect 10781 17691 10839 17697
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 13556 17737 13584 17768
rect 14550 17756 14556 17808
rect 14608 17796 14614 17808
rect 21192 17796 21220 17836
rect 22189 17833 22201 17836
rect 22235 17833 22247 17867
rect 22189 17827 22247 17833
rect 14608 17768 21220 17796
rect 14608 17756 14614 17768
rect 13541 17731 13599 17737
rect 11388 17700 12434 17728
rect 11388 17688 11394 17700
rect 8619 17632 9812 17660
rect 10505 17663 10563 17669
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 10505 17629 10517 17663
rect 10551 17629 10563 17663
rect 12406 17660 12434 17700
rect 13541 17697 13553 17731
rect 13587 17697 13599 17731
rect 15930 17728 15936 17740
rect 13541 17691 13599 17697
rect 14660 17700 15936 17728
rect 13262 17660 13268 17672
rect 12406 17632 13268 17660
rect 10505 17623 10563 17629
rect 6748 17564 8432 17592
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 6822 17524 6828 17536
rect 4571 17496 6828 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 7469 17527 7527 17533
rect 7469 17524 7481 17527
rect 6972 17496 7481 17524
rect 6972 17484 6978 17496
rect 7469 17493 7481 17496
rect 7515 17493 7527 17527
rect 8404 17524 8432 17564
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 9493 17595 9551 17601
rect 9493 17592 9505 17595
rect 8536 17564 9505 17592
rect 8536 17552 8542 17564
rect 9493 17561 9505 17564
rect 9539 17561 9551 17595
rect 9493 17555 9551 17561
rect 9582 17552 9588 17604
rect 9640 17592 9646 17604
rect 10137 17595 10195 17601
rect 10137 17592 10149 17595
rect 9640 17564 10149 17592
rect 9640 17552 9646 17564
rect 10137 17561 10149 17564
rect 10183 17561 10195 17595
rect 10520 17592 10548 17623
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 14090 17660 14096 17672
rect 13403 17632 14096 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14660 17669 14688 17700
rect 15930 17688 15936 17700
rect 15988 17688 15994 17740
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17728 17463 17731
rect 17586 17728 17592 17740
rect 17451 17700 17592 17728
rect 17451 17697 17463 17700
rect 17405 17691 17463 17697
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 18598 17688 18604 17740
rect 18656 17688 18662 17740
rect 19058 17688 19064 17740
rect 19116 17728 19122 17740
rect 20073 17731 20131 17737
rect 20073 17728 20085 17731
rect 19116 17700 20085 17728
rect 19116 17688 19122 17700
rect 20073 17697 20085 17700
rect 20119 17728 20131 17731
rect 23566 17728 23572 17740
rect 20119 17700 23572 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24854 17728 24860 17740
rect 23891 17700 24860 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17697 25191 17731
rect 25133 17691 25191 17697
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 15746 17620 15752 17672
rect 15804 17660 15810 17672
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15804 17632 16129 17660
rect 15804 17620 15810 17632
rect 16117 17629 16129 17632
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 17770 17660 17776 17672
rect 17175 17632 17776 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 17770 17620 17776 17632
rect 17828 17660 17834 17672
rect 18322 17660 18328 17672
rect 17828 17632 18328 17660
rect 17828 17620 17834 17632
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 18690 17660 18696 17672
rect 18555 17632 18696 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19518 17620 19524 17672
rect 19576 17620 19582 17672
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17660 20499 17663
rect 21450 17660 21456 17672
rect 20487 17632 21456 17660
rect 20487 17629 20499 17632
rect 20441 17623 20499 17629
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17660 21603 17663
rect 22554 17660 22560 17672
rect 21591 17632 22560 17660
rect 21591 17629 21603 17632
rect 21545 17623 21603 17629
rect 22554 17620 22560 17632
rect 22612 17620 22618 17672
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 23584 17660 23612 17688
rect 25148 17660 25176 17691
rect 23584 17632 25176 17660
rect 10520 17564 10640 17592
rect 10137 17555 10195 17561
rect 9674 17524 9680 17536
rect 8404 17496 9680 17524
rect 7469 17487 7527 17493
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 10612 17524 10640 17564
rect 11238 17552 11244 17604
rect 11296 17552 11302 17604
rect 12529 17595 12587 17601
rect 12529 17561 12541 17595
rect 12575 17561 12587 17595
rect 12529 17555 12587 17561
rect 11698 17524 11704 17536
rect 10612 17496 11704 17524
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 12544 17524 12572 17555
rect 13446 17552 13452 17604
rect 13504 17592 13510 17604
rect 13906 17592 13912 17604
rect 13504 17564 13912 17592
rect 13504 17552 13510 17564
rect 13906 17552 13912 17564
rect 13964 17592 13970 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 13964 17564 14289 17592
rect 13964 17552 13970 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 14277 17555 14335 17561
rect 16301 17595 16359 17601
rect 16301 17561 16313 17595
rect 16347 17592 16359 17595
rect 16390 17592 16396 17604
rect 16347 17564 16396 17592
rect 16347 17561 16359 17564
rect 16301 17555 16359 17561
rect 16390 17552 16396 17564
rect 16448 17552 16454 17604
rect 15470 17524 15476 17536
rect 12124 17496 15476 17524
rect 12124 17484 12130 17496
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 16758 17484 16764 17536
rect 16816 17484 16822 17536
rect 16942 17484 16948 17536
rect 17000 17524 17006 17536
rect 17126 17524 17132 17536
rect 17000 17496 17132 17524
rect 17000 17484 17006 17496
rect 17126 17484 17132 17496
rect 17184 17524 17190 17536
rect 17221 17527 17279 17533
rect 17221 17524 17233 17527
rect 17184 17496 17233 17524
rect 17184 17484 17190 17496
rect 17221 17493 17233 17496
rect 17267 17524 17279 17527
rect 17310 17524 17316 17536
rect 17267 17496 17316 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 18012 17496 18061 17524
rect 18012 17484 18018 17496
rect 18049 17493 18061 17496
rect 18095 17493 18107 17527
rect 18049 17487 18107 17493
rect 18322 17484 18328 17536
rect 18380 17524 18386 17536
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 18380 17496 18429 17524
rect 18380 17484 18386 17496
rect 18417 17493 18429 17496
rect 18463 17493 18475 17527
rect 18417 17487 18475 17493
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 19613 17527 19671 17533
rect 19613 17524 19625 17527
rect 19116 17496 19625 17524
rect 19116 17484 19122 17496
rect 19613 17493 19625 17496
rect 19659 17493 19671 17527
rect 19613 17487 19671 17493
rect 24578 17484 24584 17536
rect 24636 17484 24642 17536
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 5350 17320 5356 17332
rect 3620 17292 5356 17320
rect 3620 17193 3648 17292
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 5994 17280 6000 17332
rect 6052 17280 6058 17332
rect 6270 17280 6276 17332
rect 6328 17320 6334 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 6328 17292 6377 17320
rect 6328 17280 6334 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 8665 17323 8723 17329
rect 8665 17289 8677 17323
rect 8711 17320 8723 17323
rect 8938 17320 8944 17332
rect 8711 17292 8944 17320
rect 8711 17289 8723 17292
rect 8665 17283 8723 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9950 17280 9956 17332
rect 10008 17280 10014 17332
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 10100 17292 10425 17320
rect 10100 17280 10106 17292
rect 10413 17289 10425 17292
rect 10459 17289 10471 17323
rect 10413 17283 10471 17289
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 12802 17320 12808 17332
rect 10919 17292 12808 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 13817 17323 13875 17329
rect 13817 17289 13829 17323
rect 13863 17320 13875 17323
rect 15562 17320 15568 17332
rect 13863 17292 15568 17320
rect 13863 17289 13875 17292
rect 13817 17283 13875 17289
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 15988 17292 18889 17320
rect 15988 17280 15994 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 18877 17283 18935 17289
rect 20349 17323 20407 17329
rect 20349 17289 20361 17323
rect 20395 17320 20407 17323
rect 20395 17292 22876 17320
rect 20395 17289 20407 17292
rect 20349 17283 20407 17289
rect 6288 17252 6316 17280
rect 4080 17224 6316 17252
rect 4080 17193 4108 17224
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 9033 17255 9091 17261
rect 6880 17224 8984 17252
rect 6880 17212 6886 17224
rect 8956 17196 8984 17224
rect 9033 17221 9045 17255
rect 9079 17252 9091 17255
rect 9122 17252 9128 17264
rect 9079 17224 9128 17252
rect 9079 17221 9091 17224
rect 9033 17215 9091 17221
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 9858 17252 9864 17264
rect 9232 17224 9864 17252
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17153 3663 17187
rect 3605 17147 3663 17153
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 5350 17144 5356 17196
rect 5408 17144 5414 17196
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 5960 17156 7573 17184
rect 5960 17144 5966 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 8938 17144 8944 17196
rect 8996 17144 9002 17196
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4430 17116 4436 17128
rect 4387 17088 4436 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 2792 17048 2820 17079
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 6549 17119 6607 17125
rect 6549 17116 6561 17119
rect 5868 17088 6561 17116
rect 5868 17076 5874 17088
rect 6549 17085 6561 17088
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17116 6975 17119
rect 8294 17116 8300 17128
rect 6963 17088 8300 17116
rect 6963 17085 6975 17088
rect 6917 17079 6975 17085
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 9125 17119 9183 17125
rect 8864 17088 9076 17116
rect 8864 17048 8892 17088
rect 2792 17020 8892 17048
rect 9048 17048 9076 17088
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 9232 17116 9260 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 10137 17255 10195 17261
rect 10137 17221 10149 17255
rect 10183 17252 10195 17255
rect 11330 17252 11336 17264
rect 10183 17224 11336 17252
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 11698 17212 11704 17264
rect 11756 17252 11762 17264
rect 12526 17252 12532 17264
rect 11756 17224 12532 17252
rect 11756 17212 11762 17224
rect 12526 17212 12532 17224
rect 12584 17252 12590 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 12584 17224 13185 17252
rect 12584 17212 12590 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 13173 17215 13231 17221
rect 14185 17255 14243 17261
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 16117 17255 16175 17261
rect 16117 17252 16129 17255
rect 14231 17224 16129 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 16117 17221 16129 17224
rect 16163 17221 16175 17255
rect 22186 17252 22192 17264
rect 16117 17215 16175 17221
rect 17236 17224 19334 17252
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 10827 17156 11928 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 9171 17088 9260 17116
rect 9309 17119 9367 17125
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 9398 17116 9404 17128
rect 9355 17088 9404 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10376 17088 10977 17116
rect 10376 17076 10382 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17085 11851 17119
rect 11900 17116 11928 17156
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12032 17156 12449 17184
rect 12032 17144 12038 17156
rect 12437 17153 12449 17156
rect 12483 17184 12495 17187
rect 13906 17184 13912 17196
rect 12483 17156 13912 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 17236 17184 17264 17224
rect 15120 17156 17264 17184
rect 17405 17187 17463 17193
rect 12618 17116 12624 17128
rect 11900 17088 12624 17116
rect 11793 17079 11851 17085
rect 11514 17048 11520 17060
rect 9048 17020 11520 17048
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 2682 16940 2688 16992
rect 2740 16980 2746 16992
rect 3421 16983 3479 16989
rect 3421 16980 3433 16983
rect 2740 16952 3433 16980
rect 2740 16940 2746 16952
rect 3421 16949 3433 16952
rect 3467 16949 3479 16983
rect 3421 16943 3479 16949
rect 3602 16940 3608 16992
rect 3660 16980 3666 16992
rect 6730 16980 6736 16992
rect 3660 16952 6736 16980
rect 3660 16940 3666 16952
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 8202 16940 8208 16992
rect 8260 16940 8266 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 9674 16980 9680 16992
rect 8352 16952 9680 16980
rect 8352 16940 8358 16952
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 11808 16980 11836 17079
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17116 14335 17119
rect 14366 17116 14372 17128
rect 14323 17088 14372 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 14461 17119 14519 17125
rect 14461 17085 14473 17119
rect 14507 17116 14519 17119
rect 14734 17116 14740 17128
rect 14507 17088 14740 17116
rect 14507 17085 14519 17088
rect 14461 17079 14519 17085
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 11882 17008 11888 17060
rect 11940 17048 11946 17060
rect 15120 17048 15148 17156
rect 17405 17153 17417 17187
rect 17451 17184 17463 17187
rect 17770 17184 17776 17196
rect 17451 17156 17776 17184
rect 17451 17153 17463 17156
rect 17405 17147 17463 17153
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 17494 17076 17500 17128
rect 17552 17076 17558 17128
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17116 17739 17119
rect 17862 17116 17868 17128
rect 17727 17088 17868 17116
rect 17727 17085 17739 17088
rect 17681 17079 17739 17085
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 11940 17020 15148 17048
rect 15657 17051 15715 17057
rect 11940 17008 11946 17020
rect 15657 17017 15669 17051
rect 15703 17048 15715 17051
rect 18248 17048 18276 17147
rect 19306 17116 19334 17224
rect 19720 17224 22192 17252
rect 19720 17193 19748 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22848 17252 22876 17292
rect 22922 17280 22928 17332
rect 22980 17280 22986 17332
rect 23569 17323 23627 17329
rect 23569 17289 23581 17323
rect 23615 17320 23627 17323
rect 23842 17320 23848 17332
rect 23615 17292 23848 17320
rect 23615 17289 23627 17292
rect 23569 17283 23627 17289
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 24302 17252 24308 17264
rect 22848 17224 24308 17252
rect 24302 17212 24308 17224
rect 24360 17212 24366 17264
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 21266 17184 21272 17196
rect 20855 17156 21272 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21450 17144 21456 17196
rect 21508 17144 21514 17196
rect 22002 17144 22008 17196
rect 22060 17184 22066 17196
rect 22097 17187 22155 17193
rect 22097 17184 22109 17187
rect 22060 17156 22109 17184
rect 22060 17144 22066 17156
rect 22097 17153 22109 17156
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 19306 17088 21925 17116
rect 21913 17085 21925 17088
rect 21959 17116 21971 17119
rect 22848 17116 22876 17147
rect 23382 17144 23388 17196
rect 23440 17184 23446 17196
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23440 17156 23949 17184
rect 23440 17144 23446 17156
rect 23937 17153 23949 17156
rect 23983 17184 23995 17187
rect 24026 17184 24032 17196
rect 23983 17156 24032 17184
rect 23983 17153 23995 17156
rect 23937 17147 23995 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 25130 17184 25136 17196
rect 24688 17156 25136 17184
rect 21959 17088 22876 17116
rect 23109 17119 23167 17125
rect 21959 17085 21971 17088
rect 21913 17079 21971 17085
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 23474 17116 23480 17128
rect 23155 17088 23480 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 23474 17076 23480 17088
rect 23532 17116 23538 17128
rect 24688 17116 24716 17156
rect 25130 17144 25136 17156
rect 25188 17144 25194 17196
rect 23532 17088 24716 17116
rect 23532 17076 23538 17088
rect 24762 17076 24768 17128
rect 24820 17076 24826 17128
rect 15703 17020 18276 17048
rect 15703 17017 15715 17020
rect 15657 17011 15715 17017
rect 18414 17008 18420 17060
rect 18472 17048 18478 17060
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 18472 17020 19349 17048
rect 18472 17008 18478 17020
rect 19337 17017 19349 17020
rect 19383 17017 19395 17051
rect 19337 17011 19395 17017
rect 22462 17008 22468 17060
rect 22520 17008 22526 17060
rect 14642 16980 14648 16992
rect 11808 16952 14648 16980
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 14792 16952 16681 16980
rect 14792 16940 14798 16952
rect 16669 16949 16681 16952
rect 16715 16980 16727 16983
rect 16942 16980 16948 16992
rect 16715 16952 16948 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17037 16983 17095 16989
rect 17037 16949 17049 16983
rect 17083 16980 17095 16983
rect 17402 16980 17408 16992
rect 17083 16952 17408 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 19153 16983 19211 16989
rect 19153 16980 19165 16983
rect 17552 16952 19165 16980
rect 17552 16940 17558 16952
rect 19153 16949 19165 16952
rect 19199 16949 19211 16983
rect 19153 16943 19211 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5626 16736 5632 16788
rect 5684 16776 5690 16788
rect 5684 16748 7696 16776
rect 5684 16736 5690 16748
rect 5534 16708 5540 16720
rect 3988 16680 5540 16708
rect 3988 16649 4016 16680
rect 5534 16668 5540 16680
rect 5592 16668 5598 16720
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 7668 16708 7696 16748
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8113 16779 8171 16785
rect 8113 16776 8125 16779
rect 7800 16748 8125 16776
rect 7800 16736 7806 16748
rect 8113 16745 8125 16748
rect 8159 16745 8171 16779
rect 8113 16739 8171 16745
rect 8220 16748 11836 16776
rect 8220 16708 8248 16748
rect 6052 16680 6500 16708
rect 7668 16680 8248 16708
rect 6052 16668 6058 16680
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 4338 16640 4344 16652
rect 4295 16612 4344 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 6472 16640 6500 16680
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 8352 16680 8677 16708
rect 8352 16668 8358 16680
rect 8665 16677 8677 16680
rect 8711 16677 8723 16711
rect 11054 16708 11060 16720
rect 8665 16671 8723 16677
rect 8772 16680 11060 16708
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6472 16612 6653 16640
rect 6641 16609 6653 16612
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 6730 16600 6736 16652
rect 6788 16640 6794 16652
rect 8772 16640 8800 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 11808 16708 11836 16748
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 13964 16748 14197 16776
rect 13964 16736 13970 16748
rect 14185 16745 14197 16748
rect 14231 16776 14243 16779
rect 17218 16776 17224 16788
rect 14231 16748 17224 16776
rect 14231 16745 14243 16748
rect 14185 16739 14243 16745
rect 17218 16736 17224 16748
rect 17276 16776 17282 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 17276 16748 17417 16776
rect 17276 16736 17282 16748
rect 17405 16745 17417 16748
rect 17451 16776 17463 16779
rect 19337 16779 19395 16785
rect 19337 16776 19349 16779
rect 17451 16748 19349 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 19337 16745 19349 16748
rect 19383 16776 19395 16779
rect 19702 16776 19708 16788
rect 19383 16748 19708 16776
rect 19383 16745 19395 16748
rect 19337 16739 19395 16745
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20806 16736 20812 16788
rect 20864 16776 20870 16788
rect 20993 16779 21051 16785
rect 20993 16776 21005 16779
rect 20864 16748 21005 16776
rect 20864 16736 20870 16748
rect 20993 16745 21005 16748
rect 21039 16745 21051 16779
rect 20993 16739 21051 16745
rect 22186 16736 22192 16788
rect 22244 16736 22250 16788
rect 11808 16680 12020 16708
rect 6788 16612 8432 16640
rect 6788 16600 6794 16612
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16541 5319 16575
rect 5261 16535 5319 16541
rect 5276 16504 5304 16535
rect 5902 16532 5908 16584
rect 5960 16532 5966 16584
rect 6362 16532 6368 16584
rect 6420 16532 6426 16584
rect 8404 16572 8432 16612
rect 8588 16612 8800 16640
rect 8588 16572 8616 16612
rect 9214 16600 9220 16652
rect 9272 16640 9278 16652
rect 9585 16643 9643 16649
rect 9585 16640 9597 16643
rect 9272 16612 9597 16640
rect 9272 16600 9278 16612
rect 9585 16609 9597 16612
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 8404 16544 8616 16572
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 9692 16572 9720 16603
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 11204 16612 11253 16640
rect 11204 16600 11210 16612
rect 11241 16609 11253 16612
rect 11287 16609 11299 16643
rect 11992 16640 12020 16680
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12124 16680 13308 16708
rect 12124 16668 12130 16680
rect 13280 16649 13308 16680
rect 13354 16668 13360 16720
rect 13412 16708 13418 16720
rect 14550 16708 14556 16720
rect 13412 16680 14556 16708
rect 13412 16668 13418 16680
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 16022 16668 16028 16720
rect 16080 16708 16086 16720
rect 16393 16711 16451 16717
rect 16393 16708 16405 16711
rect 16080 16680 16405 16708
rect 16080 16668 16086 16680
rect 16393 16677 16405 16680
rect 16439 16677 16451 16711
rect 16393 16671 16451 16677
rect 17129 16711 17187 16717
rect 17129 16677 17141 16711
rect 17175 16708 17187 16711
rect 24670 16708 24676 16720
rect 17175 16680 18644 16708
rect 17175 16677 17187 16680
rect 17129 16671 17187 16677
rect 13265 16643 13323 16649
rect 11992 16612 13216 16640
rect 11241 16603 11299 16609
rect 9548 16544 9720 16572
rect 10505 16575 10563 16581
rect 9548 16532 9554 16544
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 10551 16544 11805 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 11793 16541 11805 16544
rect 11839 16572 11851 16575
rect 11974 16572 11980 16584
rect 11839 16544 11980 16572
rect 11839 16541 11851 16544
rect 11793 16535 11851 16541
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 13188 16572 13216 16612
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 13998 16600 14004 16652
rect 14056 16640 14062 16652
rect 14182 16640 14188 16652
rect 14056 16612 14188 16640
rect 14056 16600 14062 16612
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16640 14703 16643
rect 16298 16640 16304 16652
rect 14691 16612 16304 16640
rect 14691 16609 14703 16612
rect 14645 16603 14703 16609
rect 16298 16600 16304 16612
rect 16356 16640 16362 16652
rect 16850 16640 16856 16652
rect 16356 16612 16856 16640
rect 16356 16600 16362 16612
rect 16850 16600 16856 16612
rect 16908 16640 16914 16652
rect 18414 16640 18420 16652
rect 16908 16612 18420 16640
rect 16908 16600 16914 16612
rect 18414 16600 18420 16612
rect 18472 16640 18478 16652
rect 18509 16643 18567 16649
rect 18509 16640 18521 16643
rect 18472 16612 18521 16640
rect 18472 16600 18478 16612
rect 18509 16609 18521 16612
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 14274 16572 14280 16584
rect 13188 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 16054 16544 17172 16572
rect 6914 16504 6920 16516
rect 5276 16476 6920 16504
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 8570 16504 8576 16516
rect 7866 16476 8576 16504
rect 8570 16464 8576 16476
rect 8628 16464 8634 16516
rect 9674 16464 9680 16516
rect 9732 16504 9738 16516
rect 14826 16504 14832 16516
rect 9732 16476 14832 16504
rect 9732 16464 9738 16476
rect 14826 16464 14832 16476
rect 14884 16464 14890 16516
rect 14921 16507 14979 16513
rect 14921 16473 14933 16507
rect 14967 16504 14979 16507
rect 15194 16504 15200 16516
rect 14967 16476 15200 16504
rect 14967 16473 14979 16476
rect 14921 16467 14979 16473
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 16945 16507 17003 16513
rect 16945 16473 16957 16507
rect 16991 16473 17003 16507
rect 17144 16504 17172 16544
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 17773 16575 17831 16581
rect 17773 16572 17785 16575
rect 17276 16544 17785 16572
rect 17276 16532 17282 16544
rect 17773 16541 17785 16544
rect 17819 16541 17831 16575
rect 18616 16572 18644 16680
rect 18984 16680 24676 16708
rect 18690 16600 18696 16652
rect 18748 16640 18754 16652
rect 18984 16649 19012 16680
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18748 16612 18981 16640
rect 18748 16600 18754 16612
rect 18969 16609 18981 16612
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 20622 16640 20628 16652
rect 20579 16612 20628 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 18616 16544 19288 16572
rect 17773 16535 17831 16541
rect 18874 16504 18880 16516
rect 17144 16476 18880 16504
rect 16945 16467 17003 16473
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 7926 16436 7932 16448
rect 3283 16408 7932 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 8478 16396 8484 16448
rect 8536 16396 8542 16448
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 9125 16439 9183 16445
rect 9125 16436 9137 16439
rect 8904 16408 9137 16436
rect 8904 16396 8910 16408
rect 9125 16405 9137 16408
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 9493 16439 9551 16445
rect 9493 16405 9505 16439
rect 9539 16436 9551 16439
rect 10042 16436 10048 16448
rect 9539 16408 10048 16436
rect 9539 16405 9551 16408
rect 9493 16399 9551 16405
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10134 16396 10140 16448
rect 10192 16396 10198 16448
rect 11514 16396 11520 16448
rect 11572 16436 11578 16448
rect 12069 16439 12127 16445
rect 12069 16436 12081 16439
rect 11572 16408 12081 16436
rect 11572 16396 11578 16408
rect 12069 16405 12081 16408
rect 12115 16405 12127 16439
rect 12069 16399 12127 16405
rect 12710 16396 12716 16448
rect 12768 16396 12774 16448
rect 13078 16396 13084 16448
rect 13136 16396 13142 16448
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 13354 16436 13360 16448
rect 13219 16408 13360 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13817 16439 13875 16445
rect 13817 16405 13829 16439
rect 13863 16436 13875 16439
rect 14366 16436 14372 16448
rect 13863 16408 14372 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 16666 16396 16672 16448
rect 16724 16436 16730 16448
rect 16960 16436 16988 16467
rect 18874 16464 18880 16476
rect 18932 16464 18938 16516
rect 19260 16504 19288 16544
rect 19702 16532 19708 16584
rect 19760 16532 19766 16584
rect 21542 16532 21548 16584
rect 21600 16532 21606 16584
rect 22649 16575 22707 16581
rect 22649 16541 22661 16575
rect 22695 16541 22707 16575
rect 24581 16575 24639 16581
rect 24581 16572 24593 16575
rect 22649 16535 22707 16541
rect 23308 16544 24593 16572
rect 22664 16504 22692 16535
rect 19260 16476 22692 16504
rect 16724 16408 16988 16436
rect 16724 16396 16730 16408
rect 17126 16396 17132 16448
rect 17184 16436 17190 16448
rect 20714 16436 20720 16448
rect 17184 16408 20720 16436
rect 17184 16396 17190 16408
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 21266 16396 21272 16448
rect 21324 16396 21330 16448
rect 21634 16396 21640 16448
rect 21692 16436 21698 16448
rect 23308 16436 23336 16544
rect 24581 16541 24593 16544
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16572 25283 16575
rect 25958 16572 25964 16584
rect 25271 16544 25964 16572
rect 25271 16541 25283 16544
rect 25225 16535 25283 16541
rect 25958 16532 25964 16544
rect 26016 16532 26022 16584
rect 23845 16507 23903 16513
rect 23845 16473 23857 16507
rect 23891 16504 23903 16507
rect 25038 16504 25044 16516
rect 23891 16476 25044 16504
rect 23891 16473 23903 16476
rect 23845 16467 23903 16473
rect 25038 16464 25044 16476
rect 25096 16464 25102 16516
rect 21692 16408 23336 16436
rect 21692 16396 21698 16408
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 4430 16232 4436 16244
rect 2096 16204 4436 16232
rect 2096 16192 2102 16204
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 5592 16204 6469 16232
rect 5592 16192 5598 16204
rect 6457 16201 6469 16204
rect 6503 16232 6515 16235
rect 6638 16232 6644 16244
rect 6503 16204 6644 16232
rect 6503 16201 6515 16204
rect 6457 16195 6515 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 9950 16232 9956 16244
rect 7800 16204 9956 16232
rect 7800 16192 7806 16204
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10686 16232 10692 16244
rect 10459 16204 10692 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 10919 16204 13921 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 13909 16195 13967 16201
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14323 16204 14780 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 3786 16124 3792 16176
rect 3844 16164 3850 16176
rect 4065 16167 4123 16173
rect 4065 16164 4077 16167
rect 3844 16136 4077 16164
rect 3844 16124 3850 16136
rect 4065 16133 4077 16136
rect 4111 16133 4123 16167
rect 4065 16127 4123 16133
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 8110 16164 8116 16176
rect 4295 16136 8116 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 8205 16167 8263 16173
rect 8205 16133 8217 16167
rect 8251 16164 8263 16167
rect 8294 16164 8300 16176
rect 8251 16136 8300 16164
rect 8251 16133 8263 16136
rect 8205 16127 8263 16133
rect 8294 16124 8300 16136
rect 8352 16124 8358 16176
rect 8478 16124 8484 16176
rect 8536 16164 8542 16176
rect 8536 16136 8694 16164
rect 8536 16124 8542 16136
rect 10134 16124 10140 16176
rect 10192 16164 10198 16176
rect 10778 16164 10784 16176
rect 10192 16136 10784 16164
rect 10192 16124 10198 16136
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 12250 16164 12256 16176
rect 11112 16136 12256 16164
rect 11112 16124 11118 16136
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 13354 16164 13360 16176
rect 13202 16136 13360 16164
rect 13354 16124 13360 16136
rect 13412 16164 13418 16176
rect 13538 16164 13544 16176
rect 13412 16136 13544 16164
rect 13412 16124 13418 16136
rect 13538 16124 13544 16136
rect 13596 16124 13602 16176
rect 13998 16124 14004 16176
rect 14056 16164 14062 16176
rect 14752 16164 14780 16204
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15657 16235 15715 16241
rect 15657 16232 15669 16235
rect 14884 16204 15669 16232
rect 14884 16192 14890 16204
rect 15657 16201 15669 16204
rect 15703 16201 15715 16235
rect 15657 16195 15715 16201
rect 16206 16192 16212 16244
rect 16264 16232 16270 16244
rect 16482 16232 16488 16244
rect 16264 16204 16488 16232
rect 16264 16192 16270 16204
rect 16482 16192 16488 16204
rect 16540 16232 16546 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 16540 16204 18061 16232
rect 16540 16192 16546 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 21177 16235 21235 16241
rect 21177 16201 21189 16235
rect 21223 16232 21235 16235
rect 21358 16232 21364 16244
rect 21223 16204 21364 16232
rect 21223 16201 21235 16204
rect 21177 16195 21235 16201
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 15010 16164 15016 16176
rect 14056 16136 14504 16164
rect 14752 16136 15016 16164
rect 14056 16124 14062 16136
rect 658 16056 664 16108
rect 716 16096 722 16108
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 716 16068 3617 16096
rect 716 16056 722 16068
rect 3605 16065 3617 16068
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 4890 16056 4896 16108
rect 4948 16056 4954 16108
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 6178 16096 6184 16108
rect 5399 16068 6184 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 6178 16056 6184 16068
rect 6236 16056 6242 16108
rect 6836 16099 6894 16105
rect 6836 16065 6848 16099
rect 6882 16096 6894 16099
rect 7742 16096 7748 16108
rect 6882 16068 7748 16096
rect 6882 16065 6894 16068
rect 6836 16059 6894 16065
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7852 16068 7941 16096
rect 842 15988 848 16040
rect 900 16028 906 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 900 16000 3433 16028
rect 900 15988 906 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 6362 15988 6368 16040
rect 6420 16028 6426 16040
rect 6638 16028 6644 16040
rect 6420 16000 6644 16028
rect 6420 15988 6426 16000
rect 6638 15988 6644 16000
rect 6696 16028 6702 16040
rect 7282 16028 7288 16040
rect 6696 16000 7288 16028
rect 6696 15988 6702 16000
rect 7282 15988 7288 16000
rect 7340 16028 7346 16040
rect 7852 16028 7880 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 11514 16096 11520 16108
rect 7929 16059 7987 16065
rect 9646 16068 11520 16096
rect 9646 16028 9674 16068
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 7340 16000 7880 16028
rect 7340 15988 7346 16000
rect 7852 15972 7880 16000
rect 8036 16000 9674 16028
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 2498 15960 2504 15972
rect 1627 15932 2504 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 2498 15920 2504 15932
rect 2556 15920 2562 15972
rect 7834 15920 7840 15972
rect 7892 15920 7898 15972
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 8036 15960 8064 16000
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 9953 16031 10011 16037
rect 9953 16028 9965 16031
rect 9824 16000 9965 16028
rect 9824 15988 9830 16000
rect 9953 15997 9965 16000
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11103 16000 11652 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 7984 15932 8064 15960
rect 7984 15920 7990 15932
rect 2130 15852 2136 15904
rect 2188 15892 2194 15904
rect 2225 15895 2283 15901
rect 2225 15892 2237 15895
rect 2188 15864 2237 15892
rect 2188 15852 2194 15864
rect 2225 15861 2237 15864
rect 2271 15861 2283 15895
rect 2225 15855 2283 15861
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 4709 15895 4767 15901
rect 4709 15892 4721 15895
rect 4212 15864 4721 15892
rect 4212 15852 4218 15864
rect 4709 15861 4721 15864
rect 4755 15861 4767 15895
rect 4709 15855 4767 15861
rect 5994 15852 6000 15904
rect 6052 15852 6058 15904
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7469 15895 7527 15901
rect 7469 15892 7481 15895
rect 6972 15864 7481 15892
rect 6972 15852 6978 15864
rect 7469 15861 7481 15864
rect 7515 15861 7527 15895
rect 7469 15855 7527 15861
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 10134 15892 10140 15904
rect 8444 15864 10140 15892
rect 8444 15852 8450 15864
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 11624 15892 11652 16000
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12023 16000 14320 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 13078 15920 13084 15972
rect 13136 15960 13142 15972
rect 13814 15960 13820 15972
rect 13136 15932 13820 15960
rect 13136 15920 13142 15932
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 14292 15960 14320 16000
rect 14366 15988 14372 16040
rect 14424 15988 14430 16040
rect 14476 16037 14504 16136
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 15194 16124 15200 16176
rect 15252 16164 15258 16176
rect 17497 16167 17555 16173
rect 17497 16164 17509 16167
rect 15252 16136 17509 16164
rect 15252 16124 15258 16136
rect 17497 16133 17509 16136
rect 17543 16133 17555 16167
rect 17497 16127 17555 16133
rect 18230 16124 18236 16176
rect 18288 16164 18294 16176
rect 18782 16164 18788 16176
rect 18288 16136 18788 16164
rect 18288 16124 18294 16136
rect 18782 16124 18788 16136
rect 18840 16164 18846 16176
rect 18840 16136 19182 16164
rect 18840 16124 18846 16136
rect 20806 16124 20812 16176
rect 20864 16164 20870 16176
rect 20864 16136 22140 16164
rect 20864 16124 20870 16136
rect 16301 16099 16359 16105
rect 16301 16096 16313 16099
rect 15764 16068 16313 16096
rect 15764 16040 15792 16068
rect 16301 16065 16313 16068
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 16390 16056 16396 16108
rect 16448 16096 16454 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16448 16068 16865 16096
rect 16448 16056 16454 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 21082 16056 21088 16108
rect 21140 16056 21146 16108
rect 22112 16105 22140 16136
rect 25130 16124 25136 16176
rect 25188 16124 25194 16176
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 23934 16056 23940 16108
rect 23992 16056 23998 16108
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 15997 14519 16031
rect 14461 15991 14519 15997
rect 15212 16000 15424 16028
rect 15212 15960 15240 16000
rect 14292 15932 15240 15960
rect 15286 15920 15292 15972
rect 15344 15920 15350 15972
rect 15396 15960 15424 16000
rect 15746 15988 15752 16040
rect 15804 15988 15810 16040
rect 15838 15988 15844 16040
rect 15896 15988 15902 16040
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 18003 16000 18460 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 18432 15972 18460 16000
rect 18690 15988 18696 16040
rect 18748 15988 18754 16040
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19392 16000 20852 16028
rect 19392 15988 19398 16000
rect 15930 15960 15936 15972
rect 15396 15932 15936 15960
rect 15930 15920 15936 15932
rect 15988 15920 15994 15972
rect 16206 15920 16212 15972
rect 16264 15960 16270 15972
rect 16264 15932 18184 15960
rect 16264 15920 16270 15932
rect 11974 15892 11980 15904
rect 11624 15864 11980 15892
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 12768 15864 13461 15892
rect 12768 15852 12774 15864
rect 13449 15861 13461 15864
rect 13495 15892 13507 15895
rect 13722 15892 13728 15904
rect 13495 15864 13728 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 16850 15892 16856 15904
rect 15068 15864 16856 15892
rect 15068 15852 15074 15864
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 18156 15892 18184 15932
rect 18414 15920 18420 15972
rect 18472 15920 18478 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 19720 15932 20729 15960
rect 19720 15892 19748 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20824 15960 20852 16000
rect 21266 15988 21272 16040
rect 21324 16028 21330 16040
rect 21361 16031 21419 16037
rect 21361 16028 21373 16031
rect 21324 16000 21373 16028
rect 21324 15988 21330 16000
rect 21361 15997 21373 16000
rect 21407 16028 21419 16031
rect 21634 16028 21640 16040
rect 21407 16000 21640 16028
rect 21407 15997 21419 16000
rect 21361 15991 21419 15997
rect 21634 15988 21640 16000
rect 21692 15988 21698 16040
rect 23290 15988 23296 16040
rect 23348 15988 23354 16040
rect 21818 15960 21824 15972
rect 20824 15932 21824 15960
rect 20717 15923 20775 15929
rect 21818 15920 21824 15932
rect 21876 15920 21882 15972
rect 18156 15864 19748 15892
rect 20165 15895 20223 15901
rect 20165 15861 20177 15895
rect 20211 15892 20223 15895
rect 20438 15892 20444 15904
rect 20211 15864 20444 15892
rect 20211 15861 20223 15864
rect 20165 15855 20223 15861
rect 20438 15852 20444 15864
rect 20496 15892 20502 15904
rect 20806 15892 20812 15904
rect 20496 15864 20812 15892
rect 20496 15852 20502 15864
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 566 15648 572 15700
rect 624 15688 630 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 624 15660 3341 15688
rect 624 15648 630 15660
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 3329 15651 3387 15657
rect 5077 15691 5135 15697
rect 5077 15657 5089 15691
rect 5123 15688 5135 15691
rect 5350 15688 5356 15700
rect 5123 15660 5356 15688
rect 5123 15657 5135 15660
rect 5077 15651 5135 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 6178 15648 6184 15700
rect 6236 15648 6242 15700
rect 6288 15660 8432 15688
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 3418 15620 3424 15632
rect 2915 15592 3424 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 3418 15580 3424 15592
rect 3476 15580 3482 15632
rect 1949 15555 2007 15561
rect 1949 15521 1961 15555
rect 1995 15552 2007 15555
rect 3326 15552 3332 15564
rect 1995 15524 3332 15552
rect 1995 15521 2007 15524
rect 1949 15515 2007 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 750 15444 756 15496
rect 808 15484 814 15496
rect 2593 15487 2651 15493
rect 2593 15484 2605 15487
rect 808 15456 2605 15484
rect 808 15444 814 15456
rect 2593 15453 2605 15456
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 4430 15444 4436 15496
rect 4488 15444 4494 15496
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15484 5595 15487
rect 6288 15484 6316 15660
rect 8404 15629 8432 15660
rect 8754 15648 8760 15700
rect 8812 15648 8818 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 9088 15660 9137 15688
rect 9088 15648 9094 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 9548 15660 9904 15688
rect 9548 15648 9554 15660
rect 8389 15623 8447 15629
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 9398 15620 9404 15632
rect 8435 15592 9404 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 9398 15580 9404 15592
rect 9456 15580 9462 15632
rect 9769 15623 9827 15629
rect 9769 15589 9781 15623
rect 9815 15589 9827 15623
rect 9769 15583 9827 15589
rect 6638 15512 6644 15564
rect 6696 15512 6702 15564
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 9784 15552 9812 15583
rect 7340 15524 9812 15552
rect 9876 15552 9904 15660
rect 11606 15648 11612 15700
rect 11664 15688 11670 15700
rect 11793 15691 11851 15697
rect 11793 15688 11805 15691
rect 11664 15660 11805 15688
rect 11664 15648 11670 15660
rect 11793 15657 11805 15660
rect 11839 15657 11851 15691
rect 11793 15651 11851 15657
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 16206 15688 16212 15700
rect 12308 15660 16212 15688
rect 12308 15648 12314 15660
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 16408 15660 22692 15688
rect 10134 15580 10140 15632
rect 10192 15620 10198 15632
rect 11333 15623 11391 15629
rect 10192 15592 11284 15620
rect 10192 15580 10198 15592
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 9876 15524 10333 15552
rect 7340 15512 7346 15524
rect 8570 15484 8576 15496
rect 5583 15456 6316 15484
rect 8050 15456 8576 15484
rect 5583 15453 5595 15456
rect 5537 15447 5595 15453
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 8754 15444 8760 15496
rect 8812 15484 8818 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 8812 15456 9321 15484
rect 8812 15444 8818 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9876 15484 9904 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 11146 15512 11152 15564
rect 11204 15512 11210 15564
rect 9309 15447 9367 15453
rect 9416 15456 9904 15484
rect 10137 15487 10195 15493
rect 1026 15376 1032 15428
rect 1084 15416 1090 15428
rect 1673 15419 1731 15425
rect 1673 15416 1685 15419
rect 1084 15388 1685 15416
rect 1084 15376 1090 15388
rect 1673 15385 1685 15388
rect 1719 15385 1731 15419
rect 1673 15379 1731 15385
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15416 3295 15419
rect 3970 15416 3976 15428
rect 3283 15388 3976 15416
rect 3283 15385 3295 15388
rect 3237 15379 3295 15385
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 4157 15419 4215 15425
rect 4157 15385 4169 15419
rect 4203 15416 4215 15419
rect 4246 15416 4252 15428
rect 4203 15388 4252 15416
rect 4203 15385 4215 15388
rect 4157 15379 4215 15385
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 6917 15419 6975 15425
rect 6917 15385 6929 15419
rect 6963 15416 6975 15419
rect 7006 15416 7012 15428
rect 6963 15388 7012 15416
rect 6963 15385 6975 15388
rect 6917 15379 6975 15385
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 8478 15376 8484 15428
rect 8536 15416 8542 15428
rect 9416 15416 9444 15456
rect 10137 15453 10149 15487
rect 10183 15484 10195 15487
rect 11164 15484 11192 15512
rect 10183 15456 11192 15484
rect 10183 15453 10195 15456
rect 10137 15447 10195 15453
rect 8536 15388 9444 15416
rect 8536 15376 8542 15388
rect 9490 15376 9496 15428
rect 9548 15416 9554 15428
rect 11054 15416 11060 15428
rect 9548 15388 11060 15416
rect 9548 15376 9554 15388
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 11149 15419 11207 15425
rect 11149 15385 11161 15419
rect 11195 15416 11207 15419
rect 11256 15416 11284 15592
rect 11333 15589 11345 15623
rect 11379 15620 11391 15623
rect 16408 15620 16436 15660
rect 11379 15592 16436 15620
rect 11379 15589 11391 15592
rect 11333 15583 11391 15589
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 12124 15524 12357 15552
rect 12124 15512 12130 15524
rect 12345 15521 12357 15524
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 13320 15524 13400 15552
rect 13320 15512 13326 15524
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 13170 15484 13176 15496
rect 12216 15456 13176 15484
rect 12216 15444 12222 15456
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 13372 15493 13400 15524
rect 13630 15512 13636 15564
rect 13688 15512 13694 15564
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 13780 15524 14841 15552
rect 13780 15512 13786 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 16298 15512 16304 15564
rect 16356 15512 16362 15564
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 19058 15552 19064 15564
rect 16623 15524 19064 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15552 20407 15555
rect 20622 15552 20628 15564
rect 20395 15524 20628 15552
rect 20395 15521 20407 15524
rect 20349 15515 20407 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21876 15524 22109 15552
rect 21876 15512 21882 15524
rect 22097 15521 22109 15524
rect 22143 15521 22155 15555
rect 22097 15515 22155 15521
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 14642 15444 14648 15496
rect 14700 15444 14706 15496
rect 15562 15444 15568 15496
rect 15620 15444 15626 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 19242 15484 19248 15496
rect 18647 15456 19248 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 19242 15444 19248 15456
rect 19300 15484 19306 15496
rect 22664 15493 22692 15660
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19300 15456 19993 15484
rect 19300 15444 19306 15456
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 25222 15484 25228 15496
rect 24719 15456 25228 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 14737 15419 14795 15425
rect 14737 15416 14749 15419
rect 11195 15388 11284 15416
rect 13004 15388 14749 15416
rect 11195 15385 11207 15388
rect 11149 15379 11207 15385
rect 474 15308 480 15360
rect 532 15348 538 15360
rect 1489 15351 1547 15357
rect 1489 15348 1501 15351
rect 532 15320 1501 15348
rect 532 15308 538 15320
rect 1489 15317 1501 15320
rect 1535 15317 1547 15351
rect 1489 15311 1547 15317
rect 2038 15308 2044 15360
rect 2096 15308 2102 15360
rect 2222 15308 2228 15360
rect 2280 15308 2286 15360
rect 2406 15308 2412 15360
rect 2464 15308 2470 15360
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2924 15320 2973 15348
rect 2924 15308 2930 15320
rect 2961 15317 2973 15320
rect 3007 15317 3019 15351
rect 2961 15311 3019 15317
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 3694 15348 3700 15360
rect 3651 15320 3700 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 3694 15308 3700 15320
rect 3752 15308 3758 15360
rect 3878 15308 3884 15360
rect 3936 15308 3942 15360
rect 7098 15308 7104 15360
rect 7156 15348 7162 15360
rect 10134 15348 10140 15360
rect 7156 15320 10140 15348
rect 7156 15308 7162 15320
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 10229 15351 10287 15357
rect 10229 15317 10241 15351
rect 10275 15348 10287 15351
rect 10962 15348 10968 15360
rect 10275 15320 10968 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 12158 15308 12164 15360
rect 12216 15308 12222 15360
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 12526 15348 12532 15360
rect 12299 15320 12532 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 13004 15357 13032 15388
rect 14737 15385 14749 15388
rect 14783 15385 14795 15419
rect 14737 15379 14795 15385
rect 15749 15419 15807 15425
rect 15749 15385 15761 15419
rect 15795 15416 15807 15419
rect 15930 15416 15936 15428
rect 15795 15388 15936 15416
rect 15795 15385 15807 15388
rect 15749 15379 15807 15385
rect 15930 15376 15936 15388
rect 15988 15376 15994 15428
rect 18230 15416 18236 15428
rect 17802 15388 18236 15416
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 18782 15376 18788 15428
rect 18840 15376 18846 15428
rect 19518 15376 19524 15428
rect 19576 15376 19582 15428
rect 19702 15376 19708 15428
rect 19760 15376 19766 15428
rect 19886 15376 19892 15428
rect 19944 15416 19950 15428
rect 20625 15419 20683 15425
rect 20625 15416 20637 15419
rect 19944 15388 20637 15416
rect 19944 15376 19950 15388
rect 20625 15385 20637 15388
rect 20671 15385 20683 15419
rect 23845 15419 23903 15425
rect 20625 15379 20683 15385
rect 21008 15388 21114 15416
rect 21008 15360 21036 15388
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 25038 15416 25044 15428
rect 23891 15388 25044 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 25038 15376 25044 15388
rect 25096 15376 25102 15428
rect 12989 15351 13047 15357
rect 12989 15317 13001 15351
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 13449 15351 13507 15357
rect 13449 15317 13461 15351
rect 13495 15348 13507 15351
rect 13630 15348 13636 15360
rect 13495 15320 13636 15348
rect 13495 15317 13507 15320
rect 13449 15311 13507 15317
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 16022 15348 16028 15360
rect 15068 15320 16028 15348
rect 15068 15308 15074 15320
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17586 15348 17592 15360
rect 16908 15320 17592 15348
rect 16908 15308 16914 15320
rect 17586 15308 17592 15320
rect 17644 15348 17650 15360
rect 18049 15351 18107 15357
rect 18049 15348 18061 15351
rect 17644 15320 18061 15348
rect 17644 15308 17650 15320
rect 18049 15317 18061 15320
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 20990 15348 20996 15360
rect 20128 15320 20996 15348
rect 20128 15308 20134 15320
rect 20990 15308 20996 15320
rect 21048 15308 21054 15360
rect 25222 15308 25228 15360
rect 25280 15348 25286 15360
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 25280 15320 25329 15348
rect 25280 15308 25286 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 25317 15311 25375 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 4488 15116 4905 15144
rect 4488 15104 4494 15116
rect 4893 15113 4905 15116
rect 4939 15113 4951 15147
rect 4893 15107 4951 15113
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 8938 15144 8944 15156
rect 5500 15116 8944 15144
rect 5500 15104 5506 15116
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 9582 15144 9588 15156
rect 9364 15116 9588 15144
rect 9364 15104 9370 15116
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 14458 15144 14464 15156
rect 14231 15116 14464 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15381 15147 15439 15153
rect 15381 15113 15393 15147
rect 15427 15144 15439 15147
rect 15562 15144 15568 15156
rect 15427 15116 15568 15144
rect 15427 15113 15439 15116
rect 15381 15107 15439 15113
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 16390 15144 16396 15156
rect 16347 15116 16396 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 16853 15147 16911 15153
rect 16853 15113 16865 15147
rect 16899 15144 16911 15147
rect 18322 15144 18328 15156
rect 16899 15116 18328 15144
rect 16899 15113 16911 15116
rect 16853 15107 16911 15113
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 20622 15144 20628 15156
rect 19352 15116 20628 15144
rect 8386 15076 8392 15088
rect 4264 15048 8392 15076
rect 3234 14968 3240 15020
rect 3292 15008 3298 15020
rect 3878 15008 3884 15020
rect 3292 14980 3884 15008
rect 3292 14968 3298 14980
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4264 15017 4292 15048
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 8628 15048 8786 15076
rect 8628 15036 8634 15048
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10045 15079 10103 15085
rect 10045 15076 10057 15079
rect 10008 15048 10057 15076
rect 10008 15036 10014 15048
rect 10045 15045 10057 15048
rect 10091 15076 10103 15079
rect 10318 15076 10324 15088
rect 10091 15048 10324 15076
rect 10091 15045 10103 15048
rect 10045 15039 10103 15045
rect 10318 15036 10324 15048
rect 10376 15036 10382 15088
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 17221 15079 17279 15085
rect 17221 15076 17233 15079
rect 11112 15048 17233 15076
rect 11112 15036 11118 15048
rect 17221 15045 17233 15048
rect 17267 15045 17279 15079
rect 17221 15039 17279 15045
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 15008 5411 15011
rect 5994 15008 6000 15020
rect 5399 14980 6000 15008
rect 5399 14977 5411 14980
rect 5353 14971 5411 14977
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 6914 14968 6920 15020
rect 6972 14968 6978 15020
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 8021 15011 8079 15017
rect 8021 15008 8033 15011
rect 7892 14980 8033 15008
rect 7892 14968 7898 14980
rect 8021 14977 8033 14980
rect 8067 14977 8079 15011
rect 8021 14971 8079 14977
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 9640 14980 10517 15008
rect 9640 14968 9646 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11422 15008 11428 15020
rect 11195 14980 11428 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 12710 15008 12716 15020
rect 11747 14980 12716 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 15008 12863 15011
rect 12851 14980 13492 15008
rect 12851 14977 12863 14980
rect 12805 14971 12863 14977
rect 1210 14900 1216 14952
rect 1268 14940 1274 14952
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1268 14912 1961 14940
rect 1268 14900 1274 14912
rect 1949 14909 1961 14912
rect 1995 14940 2007 14943
rect 4338 14940 4344 14952
rect 1995 14912 4344 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 4338 14900 4344 14912
rect 4396 14940 4402 14952
rect 5442 14940 5448 14952
rect 4396 14912 5448 14940
rect 4396 14900 4402 14912
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 6012 14912 8309 14940
rect 934 14832 940 14884
rect 992 14872 998 14884
rect 6012 14881 6040 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 8938 14900 8944 14952
rect 8996 14940 9002 14952
rect 13464 14940 13492 14980
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 15286 15008 15292 15020
rect 14599 14980 15292 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 16574 15008 16580 15020
rect 15703 14980 16580 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 17865 15011 17923 15017
rect 17865 15008 17877 15011
rect 17328 14980 17877 15008
rect 13906 14940 13912 14952
rect 8996 14912 13400 14940
rect 13464 14912 13912 14940
rect 8996 14900 9002 14912
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 992 14844 2421 14872
rect 992 14832 998 14844
rect 2409 14841 2421 14844
rect 2455 14841 2467 14875
rect 2409 14835 2467 14841
rect 5997 14875 6055 14881
rect 5997 14841 6009 14875
rect 6043 14841 6055 14875
rect 5997 14835 6055 14841
rect 6086 14832 6092 14884
rect 6144 14872 6150 14884
rect 6457 14875 6515 14881
rect 6457 14872 6469 14875
rect 6144 14844 6469 14872
rect 6144 14832 6150 14844
rect 6457 14841 6469 14844
rect 6503 14872 6515 14875
rect 6546 14872 6552 14884
rect 6503 14844 6552 14872
rect 6503 14841 6515 14844
rect 6457 14835 6515 14841
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 6822 14872 6828 14884
rect 6687 14844 6828 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 6822 14832 6828 14844
rect 6880 14872 6886 14884
rect 7742 14872 7748 14884
rect 6880 14844 7748 14872
rect 6880 14832 6886 14844
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 13372 14872 13400 14912
rect 13906 14900 13912 14912
rect 13964 14940 13970 14952
rect 14182 14940 14188 14952
rect 13964 14912 14188 14940
rect 13964 14900 13970 14912
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14642 14900 14648 14952
rect 14700 14900 14706 14952
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 15010 14940 15016 14952
rect 14875 14912 15016 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 16206 14900 16212 14952
rect 16264 14940 16270 14952
rect 17328 14949 17356 14980
rect 17865 14977 17877 14980
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 18598 15008 18604 15020
rect 18279 14980 18604 15008
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 19352 15017 19380 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20990 15104 20996 15156
rect 21048 15144 21054 15156
rect 21048 15116 22094 15144
rect 21048 15104 21054 15116
rect 20070 15036 20076 15088
rect 20128 15036 20134 15088
rect 20898 15036 20904 15088
rect 20956 15076 20962 15088
rect 21361 15079 21419 15085
rect 21361 15076 21373 15079
rect 20956 15048 21373 15076
rect 20956 15036 20962 15048
rect 21361 15045 21373 15048
rect 21407 15045 21419 15079
rect 22066 15076 22094 15116
rect 24026 15104 24032 15156
rect 24084 15104 24090 15156
rect 22370 15076 22376 15088
rect 22066 15048 22376 15076
rect 21361 15039 21419 15045
rect 22370 15036 22376 15048
rect 22428 15076 22434 15088
rect 22428 15048 22770 15076
rect 22428 15036 22434 15048
rect 19337 15011 19395 15017
rect 19337 14977 19349 15011
rect 19383 14977 19395 15011
rect 19337 14971 19395 14977
rect 24394 14968 24400 15020
rect 24452 14968 24458 15020
rect 24670 14968 24676 15020
rect 24728 14968 24734 15020
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 16264 14912 17325 14940
rect 16264 14900 16270 14912
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 17497 14943 17555 14949
rect 17497 14909 17509 14943
rect 17543 14940 17555 14943
rect 17678 14940 17684 14952
rect 17543 14912 17684 14940
rect 17543 14909 17555 14912
rect 17497 14903 17555 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 17788 14912 19625 14940
rect 15838 14872 15844 14884
rect 9324 14844 13032 14872
rect 13372 14844 15844 14872
rect 1486 14764 1492 14816
rect 1544 14764 1550 14816
rect 1670 14764 1676 14816
rect 1728 14764 1734 14816
rect 1857 14807 1915 14813
rect 1857 14773 1869 14807
rect 1903 14804 1915 14807
rect 1946 14804 1952 14816
rect 1903 14776 1952 14804
rect 1903 14773 1915 14776
rect 1857 14767 1915 14773
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 2133 14807 2191 14813
rect 2133 14804 2145 14807
rect 2096 14776 2145 14804
rect 2096 14764 2102 14776
rect 2133 14773 2145 14776
rect 2179 14773 2191 14807
rect 2133 14767 2191 14773
rect 2590 14764 2596 14816
rect 2648 14764 2654 14816
rect 2869 14807 2927 14813
rect 2869 14773 2881 14807
rect 2915 14804 2927 14807
rect 3418 14804 3424 14816
rect 2915 14776 3424 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 6270 14804 6276 14816
rect 3835 14776 6276 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 7558 14764 7564 14816
rect 7616 14764 7622 14816
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 9324 14804 9352 14844
rect 8812 14776 9352 14804
rect 8812 14764 8818 14776
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 12345 14807 12403 14813
rect 12345 14804 12357 14807
rect 11848 14776 12357 14804
rect 11848 14764 11854 14776
rect 12345 14773 12357 14776
rect 12391 14773 12403 14807
rect 13004 14804 13032 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 16114 14832 16120 14884
rect 16172 14872 16178 14884
rect 17788 14872 17816 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 22002 14940 22008 14952
rect 20680 14912 22008 14940
rect 20680 14900 20686 14912
rect 22002 14900 22008 14912
rect 22060 14900 22066 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 22112 14912 22293 14940
rect 16172 14844 17816 14872
rect 16172 14832 16178 14844
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 20898 14872 20904 14884
rect 20772 14844 20904 14872
rect 20772 14832 20778 14844
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 22112 14872 22140 14912
rect 22281 14909 22293 14912
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 21560 14844 22140 14872
rect 21560 14816 21588 14844
rect 13354 14804 13360 14816
rect 13004 14776 13360 14804
rect 12345 14767 12403 14773
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 13630 14804 13636 14816
rect 13504 14776 13636 14804
rect 13504 14764 13510 14776
rect 13630 14764 13636 14776
rect 13688 14804 13694 14816
rect 14734 14804 14740 14816
rect 13688 14776 14740 14804
rect 13688 14764 13694 14776
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18288 14776 18889 14804
rect 18288 14764 18294 14776
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 18877 14767 18935 14773
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 21085 14807 21143 14813
rect 21085 14804 21097 14807
rect 20680 14776 21097 14804
rect 20680 14764 20686 14776
rect 21085 14773 21097 14776
rect 21131 14773 21143 14807
rect 21085 14767 21143 14773
rect 21542 14764 21548 14816
rect 21600 14764 21606 14816
rect 21634 14764 21640 14816
rect 21692 14804 21698 14816
rect 23753 14807 23811 14813
rect 23753 14804 23765 14807
rect 21692 14776 23765 14804
rect 21692 14764 21698 14776
rect 23753 14773 23765 14776
rect 23799 14773 23811 14807
rect 23753 14767 23811 14773
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 4062 14600 4068 14612
rect 3936 14572 4068 14600
rect 3936 14560 3942 14572
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 6365 14603 6423 14609
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 7006 14600 7012 14612
rect 6411 14572 7012 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 10394 14603 10452 14609
rect 10394 14600 10406 14603
rect 7616 14572 10406 14600
rect 7616 14560 7622 14572
rect 10394 14569 10406 14572
rect 10440 14569 10452 14603
rect 10394 14563 10452 14569
rect 12618 14560 12624 14612
rect 12676 14560 12682 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 13228 14572 15485 14600
rect 13228 14560 13234 14572
rect 15473 14569 15485 14572
rect 15519 14600 15531 14603
rect 15562 14600 15568 14612
rect 15519 14572 15568 14600
rect 15519 14569 15531 14572
rect 15473 14563 15531 14569
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 16574 14560 16580 14612
rect 16632 14560 16638 14612
rect 20625 14603 20683 14609
rect 20625 14569 20637 14603
rect 20671 14600 20683 14603
rect 22554 14600 22560 14612
rect 20671 14572 22560 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 22554 14560 22560 14572
rect 22612 14560 22618 14612
rect 23658 14560 23664 14612
rect 23716 14600 23722 14612
rect 23937 14603 23995 14609
rect 23937 14600 23949 14603
rect 23716 14572 23949 14600
rect 23716 14560 23722 14572
rect 23937 14569 23949 14572
rect 23983 14569 23995 14603
rect 23937 14563 23995 14569
rect 2314 14492 2320 14544
rect 2372 14532 2378 14544
rect 3237 14535 3295 14541
rect 3237 14532 3249 14535
rect 2372 14504 3249 14532
rect 2372 14492 2378 14504
rect 3237 14501 3249 14504
rect 3283 14501 3295 14535
rect 3237 14495 3295 14501
rect 4430 14492 4436 14544
rect 4488 14532 4494 14544
rect 5166 14532 5172 14544
rect 4488 14504 5172 14532
rect 4488 14492 4494 14504
rect 5166 14492 5172 14504
rect 5224 14492 5230 14544
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 7374 14532 7380 14544
rect 6052 14504 7380 14532
rect 6052 14492 6058 14504
rect 7374 14492 7380 14504
rect 7432 14492 7438 14544
rect 8573 14535 8631 14541
rect 8573 14501 8585 14535
rect 8619 14532 8631 14535
rect 9582 14532 9588 14544
rect 8619 14504 9588 14532
rect 8619 14501 8631 14504
rect 8573 14495 8631 14501
rect 9582 14492 9588 14504
rect 9640 14492 9646 14544
rect 13630 14532 13636 14544
rect 13280 14504 13636 14532
rect 6914 14464 6920 14476
rect 3436 14436 6920 14464
rect 2038 14356 2044 14408
rect 2096 14356 2102 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2682 14396 2688 14408
rect 2639 14368 2688 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3436 14405 3464 14436
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7852 14436 8248 14464
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3936 14368 3985 14396
rect 3936 14356 3942 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7852 14396 7880 14436
rect 6871 14368 7880 14396
rect 7963 14399 8021 14405
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 7963 14365 7975 14399
rect 8009 14396 8021 14399
rect 8220 14396 8248 14436
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 8996 14436 9229 14464
rect 8996 14424 9002 14436
rect 9217 14433 9229 14436
rect 9263 14464 9275 14467
rect 9306 14464 9312 14476
rect 9263 14436 9312 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 9490 14424 9496 14476
rect 9548 14424 9554 14476
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 11698 14464 11704 14476
rect 10183 14436 11704 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 11974 14424 11980 14476
rect 12032 14464 12038 14476
rect 13280 14473 13308 14504
rect 13630 14492 13636 14504
rect 13688 14532 13694 14544
rect 13998 14532 14004 14544
rect 13688 14504 14004 14532
rect 13688 14492 13694 14504
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 14182 14492 14188 14544
rect 14240 14532 14246 14544
rect 14642 14532 14648 14544
rect 14240 14504 14648 14532
rect 14240 14492 14246 14504
rect 14642 14492 14648 14504
rect 14700 14492 14706 14544
rect 15746 14532 15752 14544
rect 15580 14504 15752 14532
rect 15580 14476 15608 14504
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 21726 14532 21732 14544
rect 15856 14504 21732 14532
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 12032 14436 12173 14464
rect 12032 14424 12038 14436
rect 12161 14433 12173 14436
rect 12207 14464 12219 14467
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 12207 14436 13277 14464
rect 12207 14433 12219 14436
rect 12161 14427 12219 14433
rect 13265 14433 13277 14436
rect 13311 14433 13323 14467
rect 13265 14427 13323 14433
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 13964 14436 15056 14464
rect 13964 14424 13970 14436
rect 9766 14396 9772 14408
rect 8009 14368 8156 14396
rect 8220 14368 9772 14396
rect 8009 14365 8021 14368
rect 7963 14359 8021 14365
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 4062 14328 4068 14340
rect 2823 14300 4068 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 4062 14288 4068 14300
rect 4120 14288 4126 14340
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1489 14263 1547 14269
rect 1489 14260 1501 14263
rect 1452 14232 1501 14260
rect 1452 14220 1458 14232
rect 1489 14229 1501 14232
rect 1535 14229 1547 14263
rect 1489 14223 1547 14229
rect 1854 14220 1860 14272
rect 1912 14220 1918 14272
rect 4724 14260 4752 14359
rect 5258 14288 5264 14340
rect 5316 14288 5322 14340
rect 5736 14328 5764 14359
rect 7098 14328 7104 14340
rect 5736 14300 7104 14328
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 7650 14328 7656 14340
rect 7432 14300 7656 14328
rect 7432 14288 7438 14300
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 8128 14328 8156 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 12710 14356 12716 14408
rect 12768 14396 12774 14408
rect 14182 14396 14188 14408
rect 12768 14368 14188 14396
rect 12768 14356 12774 14368
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14458 14356 14464 14408
rect 14516 14356 14522 14408
rect 15028 14396 15056 14436
rect 15562 14424 15568 14476
rect 15620 14424 15626 14476
rect 15856 14396 15884 14504
rect 21726 14492 21732 14504
rect 21784 14492 21790 14544
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 17770 14464 17776 14476
rect 16724 14436 17776 14464
rect 16724 14424 16730 14436
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 20070 14424 20076 14476
rect 20128 14424 20134 14476
rect 21269 14467 21327 14473
rect 21269 14433 21281 14467
rect 21315 14464 21327 14467
rect 21634 14464 21640 14476
rect 21315 14436 21640 14464
rect 21315 14433 21327 14436
rect 21269 14427 21327 14433
rect 21634 14424 21640 14436
rect 21692 14424 21698 14476
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 22189 14467 22247 14473
rect 22189 14464 22201 14467
rect 22060 14436 22201 14464
rect 22060 14424 22066 14436
rect 22189 14433 22201 14436
rect 22235 14433 22247 14467
rect 22189 14427 22247 14433
rect 15028 14368 15884 14396
rect 15930 14356 15936 14408
rect 15988 14356 15994 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 16908 14368 17049 14396
rect 16908 14356 16914 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 18230 14356 18236 14408
rect 18288 14356 18294 14408
rect 19518 14356 19524 14408
rect 19576 14356 19582 14408
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20956 14368 21097 14396
rect 20956 14356 20962 14368
rect 21085 14365 21097 14368
rect 21131 14396 21143 14399
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21131 14368 21833 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14396 24639 14399
rect 25130 14396 25136 14408
rect 24627 14368 25136 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 25130 14356 25136 14368
rect 25188 14356 25194 14408
rect 12066 14328 12072 14340
rect 8128 14300 10824 14328
rect 11638 14300 12072 14328
rect 6546 14260 6552 14272
rect 4724 14232 6552 14260
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 6788 14232 7481 14260
rect 6788 14220 6794 14232
rect 7469 14229 7481 14232
rect 7515 14229 7527 14263
rect 7469 14223 7527 14229
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 7800 14232 8953 14260
rect 7800 14220 7806 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 10502 14260 10508 14272
rect 9824 14232 10508 14260
rect 9824 14220 9830 14232
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 10796 14260 10824 14300
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 12989 14331 13047 14337
rect 12989 14328 13001 14331
rect 12584 14300 13001 14328
rect 12584 14288 12590 14300
rect 12989 14297 13001 14300
rect 13035 14297 13047 14331
rect 12989 14291 13047 14297
rect 13081 14331 13139 14337
rect 13081 14297 13093 14331
rect 13127 14328 13139 14331
rect 13906 14328 13912 14340
rect 13127 14300 13912 14328
rect 13127 14297 13139 14300
rect 13081 14291 13139 14297
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 14826 14288 14832 14340
rect 14884 14328 14890 14340
rect 15565 14331 15623 14337
rect 15565 14328 15577 14331
rect 14884 14300 15577 14328
rect 14884 14288 14890 14300
rect 15565 14297 15577 14300
rect 15611 14328 15623 14331
rect 16022 14328 16028 14340
rect 15611 14300 16028 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 16022 14288 16028 14300
rect 16080 14288 16086 14340
rect 17494 14288 17500 14340
rect 17552 14328 17558 14340
rect 17552 14300 21956 14328
rect 17552 14288 17558 14300
rect 11974 14260 11980 14272
rect 10796 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13504 14232 13645 14260
rect 13504 14220 13510 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14332 14232 15117 14260
rect 14332 14220 14338 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 15470 14220 15476 14272
rect 15528 14260 15534 14272
rect 16206 14260 16212 14272
rect 15528 14232 16212 14260
rect 15528 14220 15534 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 17678 14220 17684 14272
rect 17736 14220 17742 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 18877 14263 18935 14269
rect 18877 14260 18889 14263
rect 18472 14232 18889 14260
rect 18472 14220 18478 14232
rect 18877 14229 18889 14232
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 20993 14263 21051 14269
rect 20993 14260 21005 14263
rect 20956 14232 21005 14260
rect 20956 14220 20962 14232
rect 20993 14229 21005 14232
rect 21039 14229 21051 14263
rect 21928 14260 21956 14300
rect 22002 14288 22008 14340
rect 22060 14328 22066 14340
rect 22465 14331 22523 14337
rect 22465 14328 22477 14331
rect 22060 14300 22477 14328
rect 22060 14288 22066 14300
rect 22465 14297 22477 14300
rect 22511 14297 22523 14331
rect 22465 14291 22523 14297
rect 23014 14288 23020 14340
rect 23072 14288 23078 14340
rect 22186 14260 22192 14272
rect 21928 14232 22192 14260
rect 20993 14223 21051 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 25038 14220 25044 14272
rect 25096 14260 25102 14272
rect 25225 14263 25283 14269
rect 25225 14260 25237 14263
rect 25096 14232 25237 14260
rect 25096 14220 25102 14232
rect 25225 14229 25237 14232
rect 25271 14229 25283 14263
rect 25225 14223 25283 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 1762 14056 1768 14068
rect 1719 14028 1768 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 5994 14016 6000 14068
rect 6052 14016 6058 14068
rect 6457 14059 6515 14065
rect 6457 14025 6469 14059
rect 6503 14056 6515 14059
rect 6546 14056 6552 14068
rect 6503 14028 6552 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 9398 14056 9404 14068
rect 6656 14028 9404 14056
rect 4893 13991 4951 13997
rect 4893 13957 4905 13991
rect 4939 13988 4951 13991
rect 5718 13988 5724 14000
rect 4939 13960 5724 13988
rect 4939 13957 4951 13960
rect 4893 13951 4951 13957
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13920 2375 13923
rect 2774 13920 2780 13932
rect 2363 13892 2780 13920
rect 2363 13889 2375 13892
rect 2317 13883 2375 13889
rect 2774 13880 2780 13892
rect 2832 13920 2838 13932
rect 3878 13920 3884 13932
rect 2832 13892 3884 13920
rect 2832 13880 2838 13892
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 4246 13880 4252 13932
rect 4304 13880 4310 13932
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 6270 13920 6276 13932
rect 5399 13892 6276 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 6656 13920 6684 14028
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 9548 14028 9597 14056
rect 9548 14016 9554 14028
rect 9585 14025 9597 14028
rect 9631 14025 9643 14059
rect 9585 14019 9643 14025
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 10100 14028 10425 14056
rect 10100 14016 10106 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10870 14056 10876 14068
rect 10413 14019 10471 14025
rect 10796 14028 10876 14056
rect 7742 13948 7748 14000
rect 7800 13948 7806 14000
rect 10226 13988 10232 14000
rect 8312 13960 10232 13988
rect 6733 13923 6791 13929
rect 6733 13920 6745 13923
rect 6656 13892 6745 13920
rect 6733 13889 6745 13892
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2188 13824 2605 13852
rect 2188 13812 2194 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 8312 13852 8340 13960
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 10796 13988 10824 14028
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 12345 14059 12403 14065
rect 12345 14056 12357 14059
rect 12176 14028 12357 14056
rect 12176 13988 12204 14028
rect 12345 14025 12357 14028
rect 12391 14025 12403 14059
rect 12345 14019 12403 14025
rect 12805 14059 12863 14065
rect 12805 14025 12817 14059
rect 12851 14025 12863 14059
rect 12805 14019 12863 14025
rect 12820 13988 12848 14019
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 13265 14059 13323 14065
rect 13265 14025 13277 14059
rect 13311 14056 13323 14059
rect 13354 14056 13360 14068
rect 13311 14028 13360 14056
rect 13311 14025 13323 14028
rect 13265 14019 13323 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 15252 14028 16865 14056
rect 15252 14016 15258 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 17494 14056 17500 14068
rect 17267 14028 17500 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 17494 14016 17500 14028
rect 17552 14016 17558 14068
rect 17957 14059 18015 14065
rect 17957 14025 17969 14059
rect 18003 14056 18015 14059
rect 18506 14056 18512 14068
rect 18003 14028 18512 14056
rect 18003 14025 18015 14028
rect 17957 14019 18015 14025
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 19058 14016 19064 14068
rect 19116 14016 19122 14068
rect 19334 14016 19340 14068
rect 19392 14016 19398 14068
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 19484 14028 20177 14056
rect 19484 14016 19490 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 21269 14059 21327 14065
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 23934 14056 23940 14068
rect 21315 14028 23940 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 25041 14059 25099 14065
rect 25041 14025 25053 14059
rect 25087 14056 25099 14059
rect 25774 14056 25780 14068
rect 25087 14028 25780 14056
rect 25087 14025 25099 14028
rect 25041 14019 25099 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 10612 13960 10824 13988
rect 10888 13960 12204 13988
rect 12406 13960 12848 13988
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 10612 13920 10640 13960
rect 8987 13892 10640 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10744 13892 10793 13920
rect 10744 13880 10750 13892
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 3651 13824 8340 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8444 13824 8493 13852
rect 8444 13812 8450 13824
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 8754 13784 8760 13796
rect 8076 13756 8760 13784
rect 8076 13744 8082 13756
rect 8754 13744 8760 13756
rect 8812 13744 8818 13796
rect 9140 13784 9168 13812
rect 9217 13787 9275 13793
rect 9217 13784 9229 13787
rect 9140 13756 9229 13784
rect 9217 13753 9229 13756
rect 9263 13753 9275 13787
rect 9217 13747 9275 13753
rect 9582 13744 9588 13796
rect 9640 13784 9646 13796
rect 9692 13784 9720 13815
rect 9766 13812 9772 13864
rect 9824 13812 9830 13864
rect 10888 13852 10916 13960
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 11790 13920 11796 13932
rect 11747 13892 11796 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 12406 13920 12434 13960
rect 14274 13948 14280 14000
rect 14332 13948 14338 14000
rect 14826 13948 14832 14000
rect 14884 13948 14890 14000
rect 17313 13991 17371 13997
rect 17313 13988 17325 13991
rect 15580 13960 17325 13988
rect 13446 13920 13452 13932
rect 11900 13892 12434 13920
rect 13280 13892 13452 13920
rect 9876 13824 10916 13852
rect 10965 13855 11023 13861
rect 9640 13756 9720 13784
rect 9640 13744 9646 13756
rect 6996 13719 7054 13725
rect 6996 13685 7008 13719
rect 7042 13716 7054 13719
rect 8386 13716 8392 13728
rect 7042 13688 8392 13716
rect 7042 13685 7054 13688
rect 6996 13679 7054 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 8570 13676 8576 13728
rect 8628 13716 8634 13728
rect 9876 13716 9904 13824
rect 10965 13821 10977 13855
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 10226 13744 10232 13796
rect 10284 13784 10290 13796
rect 10686 13784 10692 13796
rect 10284 13756 10692 13784
rect 10284 13744 10290 13756
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 10980 13784 11008 13815
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11900 13852 11928 13892
rect 11480 13824 11928 13852
rect 11480 13812 11486 13824
rect 11974 13812 11980 13864
rect 12032 13852 12038 13864
rect 13280 13852 13308 13892
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 12032 13824 13308 13852
rect 13357 13855 13415 13861
rect 12032 13812 12038 13824
rect 13357 13821 13369 13855
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 10836 13756 11008 13784
rect 10836 13744 10842 13756
rect 12250 13744 12256 13796
rect 12308 13784 12314 13796
rect 13372 13784 13400 13815
rect 13998 13812 14004 13864
rect 14056 13812 14062 13864
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 15580 13852 15608 13960
rect 17313 13957 17325 13960
rect 17359 13957 17371 13991
rect 17313 13951 17371 13957
rect 19518 13948 19524 14000
rect 19576 13988 19582 14000
rect 20809 13991 20867 13997
rect 20809 13988 20821 13991
rect 19576 13960 20821 13988
rect 19576 13948 19582 13960
rect 20809 13957 20821 13960
rect 20855 13988 20867 13991
rect 20855 13960 21864 13988
rect 20855 13957 20867 13960
rect 20809 13951 20867 13957
rect 21836 13932 21864 13960
rect 22094 13948 22100 14000
rect 22152 13948 22158 14000
rect 23014 13988 23020 14000
rect 22848 13960 23020 13988
rect 16390 13920 16396 13932
rect 14700 13824 15608 13852
rect 15672 13892 16396 13920
rect 14700 13812 14706 13824
rect 12308 13756 13400 13784
rect 12308 13744 12314 13756
rect 15378 13744 15384 13796
rect 15436 13784 15442 13796
rect 15672 13784 15700 13892
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 17862 13920 17868 13932
rect 16500 13892 17868 13920
rect 15749 13855 15807 13861
rect 15749 13821 15761 13855
rect 15795 13821 15807 13855
rect 15749 13815 15807 13821
rect 15436 13756 15700 13784
rect 15764 13784 15792 13815
rect 16022 13812 16028 13864
rect 16080 13852 16086 13864
rect 16500 13852 16528 13892
rect 17862 13880 17868 13892
rect 17920 13920 17926 13932
rect 18049 13923 18107 13929
rect 18049 13920 18061 13923
rect 17920 13892 18061 13920
rect 17920 13880 17926 13892
rect 18049 13889 18061 13892
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18414 13880 18420 13932
rect 18472 13880 18478 13932
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 19024 13892 20085 13920
rect 19024 13880 19030 13892
rect 20073 13889 20085 13892
rect 20119 13889 20131 13923
rect 20073 13883 20131 13889
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20496 13892 21097 13920
rect 20496 13880 20502 13892
rect 21085 13889 21097 13892
rect 21131 13920 21143 13923
rect 21453 13923 21511 13929
rect 21453 13920 21465 13923
rect 21131 13892 21465 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21453 13889 21465 13892
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 21818 13880 21824 13932
rect 21876 13920 21882 13932
rect 22848 13920 22876 13960
rect 23014 13948 23020 13960
rect 23072 13948 23078 14000
rect 23842 13948 23848 14000
rect 23900 13948 23906 14000
rect 21876 13892 22876 13920
rect 21876 13880 21882 13892
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 16080 13824 16528 13852
rect 17405 13855 17463 13861
rect 16080 13812 16086 13824
rect 17405 13821 17417 13855
rect 17451 13821 17463 13855
rect 20257 13855 20315 13861
rect 20257 13852 20269 13855
rect 17405 13815 17463 13821
rect 17512 13824 19748 13852
rect 15930 13784 15936 13796
rect 15764 13756 15936 13784
rect 15436 13744 15442 13756
rect 15930 13744 15936 13756
rect 15988 13784 15994 13796
rect 17420 13784 17448 13815
rect 15988 13756 17448 13784
rect 15988 13744 15994 13756
rect 8628 13688 9904 13716
rect 8628 13676 8634 13688
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 13354 13716 13360 13728
rect 10008 13688 13360 13716
rect 10008 13676 10014 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13446 13676 13452 13728
rect 13504 13716 13510 13728
rect 16022 13716 16028 13728
rect 13504 13688 16028 13716
rect 13504 13676 13510 13688
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 16206 13676 16212 13728
rect 16264 13676 16270 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 17512 13716 17540 13824
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 19720 13793 19748 13824
rect 19812 13824 20269 13852
rect 19705 13787 19763 13793
rect 17644 13756 19656 13784
rect 17644 13744 17650 13756
rect 16632 13688 17540 13716
rect 19628 13716 19656 13756
rect 19705 13753 19717 13787
rect 19751 13753 19763 13787
rect 19705 13747 19763 13753
rect 19812 13716 19840 13824
rect 20257 13821 20269 13824
rect 20303 13852 20315 13855
rect 20622 13852 20628 13864
rect 20303 13824 20628 13852
rect 20303 13821 20315 13824
rect 20257 13815 20315 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 20898 13812 20904 13864
rect 20956 13812 20962 13864
rect 22830 13812 22836 13864
rect 22888 13812 22894 13864
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24544 13824 24593 13852
rect 24544 13812 24550 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 21726 13744 21732 13796
rect 21784 13784 21790 13796
rect 22281 13787 22339 13793
rect 22281 13784 22293 13787
rect 21784 13756 22293 13784
rect 21784 13744 21790 13756
rect 22281 13753 22293 13756
rect 22327 13753 22339 13787
rect 22281 13747 22339 13753
rect 25222 13744 25228 13796
rect 25280 13784 25286 13796
rect 25406 13784 25412 13796
rect 25280 13756 25412 13784
rect 25280 13744 25286 13756
rect 25406 13744 25412 13756
rect 25464 13744 25470 13796
rect 19628 13688 19840 13716
rect 16632 13676 16638 13688
rect 21266 13676 21272 13728
rect 21324 13716 21330 13728
rect 23096 13719 23154 13725
rect 23096 13716 23108 13719
rect 21324 13688 23108 13716
rect 21324 13676 21330 13688
rect 23096 13685 23108 13688
rect 23142 13716 23154 13719
rect 24854 13716 24860 13728
rect 23142 13688 24860 13716
rect 23142 13685 23154 13688
rect 23096 13679 23154 13685
rect 24854 13676 24860 13688
rect 24912 13676 24918 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 2648 13484 4077 13512
rect 2648 13472 2654 13484
rect 4065 13481 4077 13484
rect 4111 13512 4123 13515
rect 4111 13484 5764 13512
rect 4111 13481 4123 13484
rect 4065 13475 4123 13481
rect 5626 13444 5632 13456
rect 2746 13416 5632 13444
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2746 13376 2774 13416
rect 5626 13404 5632 13416
rect 5684 13404 5690 13456
rect 5736 13444 5764 13484
rect 6270 13472 6276 13524
rect 6328 13472 6334 13524
rect 7742 13512 7748 13524
rect 6380 13484 7748 13512
rect 6380 13444 6408 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 9125 13515 9183 13521
rect 7984 13484 8708 13512
rect 7984 13472 7990 13484
rect 5736 13416 6408 13444
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13444 7435 13447
rect 8680 13444 8708 13484
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9214 13512 9220 13524
rect 9171 13484 9220 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 9916 13484 10425 13512
rect 9916 13472 9922 13484
rect 10413 13481 10425 13484
rect 10459 13481 10471 13515
rect 10413 13475 10471 13481
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 12250 13512 12256 13524
rect 10560 13484 12256 13512
rect 10560 13472 10566 13484
rect 12250 13472 12256 13484
rect 12308 13512 12314 13524
rect 12308 13484 12388 13512
rect 12308 13472 12314 13484
rect 11974 13444 11980 13456
rect 7423 13416 8616 13444
rect 8680 13416 11980 13444
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 2547 13348 2774 13376
rect 3237 13379 3295 13385
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3237 13345 3249 13379
rect 3283 13376 3295 13379
rect 5534 13376 5540 13388
rect 3283 13348 5540 13376
rect 3283 13345 3295 13348
rect 3237 13339 3295 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 5902 13336 5908 13388
rect 5960 13376 5966 13388
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 5960 13348 8309 13376
rect 5960 13336 5966 13348
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13345 8447 13379
rect 8588 13376 8616 13416
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 12360 13444 12388 13484
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13722 13512 13728 13524
rect 12492 13484 12940 13512
rect 12492 13472 12498 13484
rect 12912 13444 12940 13484
rect 13280 13484 13728 13512
rect 13280 13444 13308 13484
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 14148 13484 14197 13512
rect 14148 13472 14154 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14185 13475 14243 13481
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 17589 13515 17647 13521
rect 17589 13512 17601 13515
rect 16080 13484 17601 13512
rect 16080 13472 16086 13484
rect 17589 13481 17601 13484
rect 17635 13481 17647 13515
rect 17589 13475 17647 13481
rect 18874 13472 18880 13524
rect 18932 13472 18938 13524
rect 19334 13472 19340 13524
rect 19392 13472 19398 13524
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 21082 13512 21088 13524
rect 19475 13484 21088 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22646 13512 22652 13524
rect 22143 13484 22652 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 25225 13515 25283 13521
rect 25225 13512 25237 13515
rect 24176 13484 25237 13512
rect 24176 13472 24182 13484
rect 25225 13481 25237 13484
rect 25271 13481 25283 13515
rect 25225 13475 25283 13481
rect 14829 13447 14887 13453
rect 12360 13416 12664 13444
rect 12912 13416 13308 13444
rect 13372 13416 14780 13444
rect 9306 13376 9312 13388
rect 8588 13348 9312 13376
rect 8389 13339 8447 13345
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 2314 13268 2320 13320
rect 2372 13268 2378 13320
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 4154 13308 4160 13320
rect 3099 13280 4160 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4522 13268 4528 13320
rect 4580 13268 4586 13320
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 8018 13308 8024 13320
rect 7392 13280 8024 13308
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 3789 13243 3847 13249
rect 3789 13240 3801 13243
rect 3476 13212 3801 13240
rect 3476 13200 3482 13212
rect 3789 13209 3801 13212
rect 3835 13209 3847 13243
rect 3789 13203 3847 13209
rect 5166 13200 5172 13252
rect 5224 13200 5230 13252
rect 5442 13200 5448 13252
rect 5500 13240 5506 13252
rect 7392 13240 7420 13280
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 8404 13308 8432 13339
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 9674 13336 9680 13388
rect 9732 13336 9738 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 9824 13348 10977 13376
rect 9824 13336 9830 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13376 11575 13379
rect 12066 13376 12072 13388
rect 11563 13348 12072 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 12250 13336 12256 13388
rect 12308 13336 12314 13388
rect 12342 13336 12348 13388
rect 12400 13336 12406 13388
rect 8168 13280 8432 13308
rect 8168 13268 8174 13280
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 9122 13308 9128 13320
rect 8996 13280 9128 13308
rect 8996 13268 9002 13280
rect 9122 13268 9128 13280
rect 9180 13308 9186 13320
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 9180 13280 9505 13308
rect 9180 13268 9186 13280
rect 9493 13277 9505 13280
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13308 10839 13311
rect 12434 13308 12440 13320
rect 10827 13280 12440 13308
rect 10827 13277 10839 13280
rect 10781 13271 10839 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12636 13308 12664 13416
rect 13372 13308 13400 13416
rect 13630 13336 13636 13388
rect 13688 13336 13694 13388
rect 14752 13376 14780 13416
rect 14829 13413 14841 13447
rect 14875 13444 14887 13447
rect 17034 13444 17040 13456
rect 14875 13416 17040 13444
rect 14875 13413 14887 13416
rect 14829 13407 14887 13413
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 18564 13416 22692 13444
rect 18564 13404 18570 13416
rect 15841 13379 15899 13385
rect 15841 13376 15853 13379
rect 14752 13348 15853 13376
rect 15841 13345 15853 13348
rect 15887 13376 15899 13379
rect 16022 13376 16028 13388
rect 15887 13348 16028 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16114 13336 16120 13388
rect 16172 13376 16178 13388
rect 19426 13376 19432 13388
rect 16172 13348 19432 13376
rect 16172 13336 16178 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 19518 13336 19524 13388
rect 19576 13376 19582 13388
rect 19981 13379 20039 13385
rect 19981 13376 19993 13379
rect 19576 13348 19993 13376
rect 19576 13336 19582 13348
rect 19981 13345 19993 13348
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 20680 13348 21281 13376
rect 20680 13336 20686 13348
rect 21269 13345 21281 13348
rect 21315 13345 21327 13379
rect 21269 13339 21327 13345
rect 12636 13280 13400 13308
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 15930 13308 15936 13320
rect 13495 13280 15936 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 17678 13308 17684 13320
rect 16531 13280 17684 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 17770 13268 17776 13320
rect 17828 13268 17834 13320
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 5500 13212 7420 13240
rect 5500 13200 5506 13212
rect 7466 13200 7472 13252
rect 7524 13240 7530 13252
rect 8205 13243 8263 13249
rect 7524 13212 7880 13240
rect 7524 13200 7530 13212
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13172 3663 13175
rect 3878 13172 3884 13184
rect 3651 13144 3884 13172
rect 3651 13141 3663 13144
rect 3605 13135 3663 13141
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 7742 13172 7748 13184
rect 5408 13144 7748 13172
rect 5408 13132 5414 13144
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 7852 13181 7880 13212
rect 8205 13209 8217 13243
rect 8251 13240 8263 13243
rect 8754 13240 8760 13252
rect 8251 13212 8760 13240
rect 8251 13209 8263 13212
rect 8205 13203 8263 13209
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 9631 13212 11836 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 7926 13132 7932 13184
rect 7984 13172 7990 13184
rect 8938 13172 8944 13184
rect 7984 13144 8944 13172
rect 7984 13132 7990 13144
rect 8938 13132 8944 13144
rect 8996 13172 9002 13184
rect 9766 13172 9772 13184
rect 8996 13144 9772 13172
rect 8996 13132 9002 13144
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 10870 13132 10876 13184
rect 10928 13132 10934 13184
rect 11808 13181 11836 13212
rect 12066 13200 12072 13252
rect 12124 13240 12130 13252
rect 12161 13243 12219 13249
rect 12161 13240 12173 13243
rect 12124 13212 12173 13240
rect 12124 13200 12130 13212
rect 12161 13209 12173 13212
rect 12207 13209 12219 13243
rect 12161 13203 12219 13209
rect 12820 13212 14044 13240
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13141 11851 13175
rect 11793 13135 11851 13141
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12820 13172 12848 13212
rect 12032 13144 12848 13172
rect 12032 13132 12038 13144
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 12952 13144 13001 13172
rect 12952 13132 12958 13144
rect 12989 13141 13001 13144
rect 13035 13141 13047 13175
rect 12989 13135 13047 13141
rect 13354 13132 13360 13184
rect 13412 13132 13418 13184
rect 14016 13172 14044 13212
rect 14090 13200 14096 13252
rect 14148 13240 14154 13252
rect 14645 13243 14703 13249
rect 14645 13240 14657 13243
rect 14148 13212 14657 13240
rect 14148 13200 14154 13212
rect 14645 13209 14657 13212
rect 14691 13209 14703 13243
rect 14645 13203 14703 13209
rect 15470 13200 15476 13252
rect 15528 13240 15534 13252
rect 15657 13243 15715 13249
rect 15657 13240 15669 13243
rect 15528 13212 15669 13240
rect 15528 13200 15534 13212
rect 15657 13209 15669 13212
rect 15703 13209 15715 13243
rect 18248 13240 18276 13271
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 19300 13280 19901 13308
rect 19300 13268 19306 13280
rect 19889 13277 19901 13280
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 21174 13268 21180 13320
rect 21232 13268 21238 13320
rect 21284 13308 21312 13339
rect 21284 13280 21496 13308
rect 21358 13240 21364 13252
rect 18248 13212 21364 13240
rect 15657 13203 15715 13209
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 21468 13240 21496 13280
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22664 13317 22692 13416
rect 23845 13379 23903 13385
rect 23845 13345 23857 13379
rect 23891 13376 23903 13379
rect 23934 13376 23940 13388
rect 23891 13348 23940 13376
rect 23891 13345 23903 13348
rect 23845 13339 23903 13345
rect 23934 13336 23940 13348
rect 23992 13336 23998 13388
rect 22005 13311 22063 13317
rect 22005 13308 22017 13311
rect 21968 13280 22017 13308
rect 21968 13268 21974 13280
rect 22005 13277 22017 13280
rect 22051 13277 22063 13311
rect 22005 13271 22063 13277
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13277 22707 13311
rect 22649 13271 22707 13277
rect 23750 13268 23756 13320
rect 23808 13308 23814 13320
rect 24210 13308 24216 13320
rect 23808 13280 24216 13308
rect 23808 13268 23814 13280
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 24578 13268 24584 13320
rect 24636 13268 24642 13320
rect 24486 13240 24492 13252
rect 21468 13212 24492 13240
rect 24486 13200 24492 13212
rect 24544 13200 24550 13252
rect 15102 13172 15108 13184
rect 14016 13144 15108 13172
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 15252 13144 15301 13172
rect 15252 13132 15258 13144
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 15289 13135 15347 13141
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 15562 13172 15568 13184
rect 15436 13144 15568 13172
rect 15436 13132 15442 13144
rect 15562 13132 15568 13144
rect 15620 13172 15626 13184
rect 15749 13175 15807 13181
rect 15749 13172 15761 13175
rect 15620 13144 15761 13172
rect 15620 13132 15626 13144
rect 15749 13141 15761 13144
rect 15795 13141 15807 13175
rect 15749 13135 15807 13141
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 17129 13175 17187 13181
rect 17129 13172 17141 13175
rect 16908 13144 17141 13172
rect 16908 13132 16914 13144
rect 17129 13141 17141 13144
rect 17175 13141 17187 13175
rect 17129 13135 17187 13141
rect 17862 13132 17868 13184
rect 17920 13172 17926 13184
rect 19058 13172 19064 13184
rect 17920 13144 19064 13172
rect 17920 13132 17926 13144
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19797 13175 19855 13181
rect 19797 13172 19809 13175
rect 19392 13144 19809 13172
rect 19392 13132 19398 13144
rect 19797 13141 19809 13144
rect 19843 13141 19855 13175
rect 19797 13135 19855 13141
rect 20714 13132 20720 13184
rect 20772 13132 20778 13184
rect 21082 13132 21088 13184
rect 21140 13132 21146 13184
rect 22554 13132 22560 13184
rect 22612 13172 22618 13184
rect 22922 13172 22928 13184
rect 22612 13144 22928 13172
rect 22612 13132 22618 13144
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 2593 12971 2651 12977
rect 2593 12937 2605 12971
rect 2639 12937 2651 12971
rect 2593 12931 2651 12937
rect 2133 12835 2191 12841
rect 2133 12832 2145 12835
rect 1504 12804 2145 12832
rect 1118 12588 1124 12640
rect 1176 12628 1182 12640
rect 1504 12637 1532 12804
rect 2133 12801 2145 12804
rect 2179 12801 2191 12835
rect 2133 12795 2191 12801
rect 2608 12764 2636 12931
rect 3602 12928 3608 12980
rect 3660 12968 3666 12980
rect 3878 12968 3884 12980
rect 3660 12940 3884 12968
rect 3660 12928 3666 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 4856 12940 7604 12968
rect 4856 12928 4862 12940
rect 3237 12903 3295 12909
rect 3237 12869 3249 12903
rect 3283 12900 3295 12903
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 3283 12872 7481 12900
rect 3283 12869 3295 12872
rect 3237 12863 3295 12869
rect 7469 12869 7481 12872
rect 7515 12869 7527 12903
rect 7576 12900 7604 12940
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 8662 12968 8668 12980
rect 7800 12940 8668 12968
rect 7800 12928 7806 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9398 12928 9404 12980
rect 9456 12968 9462 12980
rect 10502 12968 10508 12980
rect 9456 12940 10508 12968
rect 9456 12928 9462 12940
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12216 12940 13093 12968
rect 12216 12928 12222 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 13081 12931 13139 12937
rect 13446 12928 13452 12980
rect 13504 12928 13510 12980
rect 14182 12928 14188 12980
rect 14240 12968 14246 12980
rect 16574 12968 16580 12980
rect 14240 12940 16580 12968
rect 14240 12928 14246 12940
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 18138 12968 18144 12980
rect 17512 12940 18144 12968
rect 9766 12900 9772 12912
rect 7576 12872 9772 12900
rect 7469 12863 7527 12869
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 10134 12860 10140 12912
rect 10192 12860 10198 12912
rect 11701 12903 11759 12909
rect 11701 12869 11713 12903
rect 11747 12900 11759 12903
rect 11882 12900 11888 12912
rect 11747 12872 11888 12900
rect 11747 12869 11759 12872
rect 11701 12863 11759 12869
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 12342 12860 12348 12912
rect 12400 12900 12406 12912
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 12400 12872 12449 12900
rect 12400 12860 12406 12872
rect 12437 12869 12449 12872
rect 12483 12869 12495 12903
rect 12437 12863 12495 12869
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 15933 12903 15991 12909
rect 14424 12872 14964 12900
rect 14424 12860 14430 12872
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3786 12832 3792 12844
rect 2823 12804 3792 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 5074 12832 5080 12844
rect 4295 12804 5080 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 8297 12835 8355 12841
rect 5644 12804 7788 12832
rect 5644 12764 5672 12804
rect 2608 12736 5672 12764
rect 6822 12724 6828 12776
rect 6880 12724 6886 12776
rect 7558 12724 7564 12776
rect 7616 12724 7622 12776
rect 7650 12724 7656 12776
rect 7708 12724 7714 12776
rect 7760 12764 7788 12804
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 8570 12832 8576 12844
rect 8343 12804 8576 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 13556 12804 14749 12832
rect 8478 12764 8484 12776
rect 7760 12736 8484 12764
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 8987 12736 9689 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 11992 12764 12020 12792
rect 13556 12773 13584 12804
rect 14737 12801 14749 12804
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 9677 12727 9735 12733
rect 11072 12736 12020 12764
rect 12084 12736 13553 12764
rect 1673 12699 1731 12705
rect 1673 12665 1685 12699
rect 1719 12696 1731 12699
rect 1762 12696 1768 12708
rect 1719 12668 1768 12696
rect 1719 12665 1731 12668
rect 1673 12659 1731 12665
rect 1762 12656 1768 12668
rect 1820 12656 1826 12708
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 5442 12696 5448 12708
rect 1995 12668 5448 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 6457 12699 6515 12705
rect 6457 12696 6469 12699
rect 5684 12668 6469 12696
rect 5684 12656 5690 12668
rect 6457 12665 6469 12668
rect 6503 12696 6515 12699
rect 6503 12668 8156 12696
rect 6503 12665 6515 12668
rect 6457 12659 6515 12665
rect 1489 12631 1547 12637
rect 1489 12628 1501 12631
rect 1176 12600 1501 12628
rect 1176 12588 1182 12600
rect 1489 12597 1501 12600
rect 1535 12597 1547 12631
rect 1489 12591 1547 12597
rect 3786 12588 3792 12640
rect 3844 12588 3850 12640
rect 4893 12631 4951 12637
rect 4893 12597 4905 12631
rect 4939 12628 4951 12631
rect 5350 12628 5356 12640
rect 4939 12600 5356 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 5994 12588 6000 12640
rect 6052 12588 6058 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 6546 12628 6552 12640
rect 6420 12600 6552 12628
rect 6420 12588 6426 12600
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 6638 12588 6644 12640
rect 6696 12588 6702 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7742 12628 7748 12640
rect 7147 12600 7748 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 8128 12628 8156 12668
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 8754 12696 8760 12708
rect 8260 12668 8760 12696
rect 8260 12656 8266 12668
rect 8754 12656 8760 12668
rect 8812 12656 8818 12708
rect 11072 12628 11100 12736
rect 11698 12656 11704 12708
rect 11756 12696 11762 12708
rect 12084 12696 12112 12736
rect 13541 12733 13553 12736
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 13722 12724 13728 12776
rect 13780 12724 13786 12776
rect 14826 12724 14832 12776
rect 14884 12724 14890 12776
rect 14936 12773 14964 12872
rect 15933 12869 15945 12903
rect 15979 12900 15991 12903
rect 17512 12900 17540 12940
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 18414 12928 18420 12980
rect 18472 12968 18478 12980
rect 19242 12968 19248 12980
rect 18472 12940 19248 12968
rect 18472 12928 18478 12940
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 20622 12968 20628 12980
rect 19484 12940 20628 12968
rect 19484 12928 19490 12940
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 21910 12928 21916 12980
rect 21968 12968 21974 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 21968 12940 25237 12968
rect 21968 12928 21974 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 25225 12931 25283 12937
rect 15979 12872 17540 12900
rect 15979 12869 15991 12872
rect 15933 12863 15991 12869
rect 17862 12860 17868 12912
rect 17920 12860 17926 12912
rect 18874 12860 18880 12912
rect 18932 12900 18938 12912
rect 19058 12900 19064 12912
rect 18932 12872 19064 12900
rect 18932 12860 18938 12872
rect 19058 12860 19064 12872
rect 19116 12860 19122 12912
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19610 12900 19616 12912
rect 19392 12872 19616 12900
rect 19392 12860 19398 12872
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 19794 12860 19800 12912
rect 19852 12900 19858 12912
rect 21085 12903 21143 12909
rect 21085 12900 21097 12903
rect 19852 12872 21097 12900
rect 19852 12860 19858 12872
rect 21085 12869 21097 12872
rect 21131 12869 21143 12903
rect 21085 12863 21143 12869
rect 21637 12903 21695 12909
rect 21637 12869 21649 12903
rect 21683 12900 21695 12903
rect 22002 12900 22008 12912
rect 21683 12872 22008 12900
rect 21683 12869 21695 12872
rect 21637 12863 21695 12869
rect 22002 12860 22008 12872
rect 22060 12860 22066 12912
rect 22370 12900 22376 12912
rect 22112 12872 22376 12900
rect 22112 12844 22140 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 23290 12860 23296 12912
rect 23348 12860 23354 12912
rect 23842 12860 23848 12912
rect 23900 12860 23906 12912
rect 24578 12860 24584 12912
rect 24636 12900 24642 12912
rect 25041 12903 25099 12909
rect 25041 12900 25053 12903
rect 24636 12872 25053 12900
rect 24636 12860 24642 12872
rect 25041 12869 25053 12872
rect 25087 12869 25099 12903
rect 25041 12863 25099 12869
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16206 12832 16212 12844
rect 16071 12804 16212 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 18340 12804 20576 12832
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 16114 12724 16120 12776
rect 16172 12724 16178 12776
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 11756 12668 12112 12696
rect 11756 12656 11762 12668
rect 12158 12656 12164 12708
rect 12216 12696 12222 12708
rect 15565 12699 15623 12705
rect 15565 12696 15577 12699
rect 12216 12668 15577 12696
rect 12216 12656 12222 12668
rect 15565 12665 15577 12668
rect 15611 12665 15623 12699
rect 15565 12659 15623 12665
rect 8128 12600 11100 12628
rect 11146 12588 11152 12640
rect 11204 12588 11210 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 14182 12628 14188 12640
rect 11664 12600 14188 12628
rect 11664 12588 11670 12600
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 14369 12631 14427 12637
rect 14369 12597 14381 12631
rect 14415 12628 14427 12631
rect 14642 12628 14648 12640
rect 14415 12600 14648 12628
rect 14415 12597 14427 12600
rect 14369 12591 14427 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 16574 12628 16580 12640
rect 15160 12600 16580 12628
rect 15160 12588 15166 12600
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16868 12628 16896 12727
rect 17126 12724 17132 12776
rect 17184 12724 17190 12776
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 18340 12764 18368 12804
rect 17276 12736 18368 12764
rect 17276 12724 17282 12736
rect 20438 12724 20444 12776
rect 20496 12724 20502 12776
rect 20548 12764 20576 12804
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 24912 12804 25421 12832
rect 24912 12792 24918 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 21818 12764 21824 12776
rect 20548 12736 21824 12764
rect 21818 12724 21824 12736
rect 21876 12724 21882 12776
rect 21910 12724 21916 12776
rect 21968 12764 21974 12776
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 21968 12736 22293 12764
rect 21968 12724 21974 12736
rect 22281 12733 22293 12736
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 22646 12724 22652 12776
rect 22704 12764 22710 12776
rect 22830 12764 22836 12776
rect 22704 12736 22836 12764
rect 22704 12724 22710 12736
rect 22830 12724 22836 12736
rect 22888 12764 22894 12776
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22888 12736 23029 12764
rect 22888 12724 22894 12736
rect 23017 12733 23029 12736
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 23842 12724 23848 12776
rect 23900 12764 23906 12776
rect 24486 12764 24492 12776
rect 23900 12736 24492 12764
rect 23900 12724 23906 12736
rect 24486 12724 24492 12736
rect 24544 12724 24550 12776
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 18969 12699 19027 12705
rect 18969 12696 18981 12699
rect 18196 12668 18981 12696
rect 18196 12656 18202 12668
rect 18969 12665 18981 12668
rect 19015 12696 19027 12699
rect 19015 12668 19564 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 18506 12628 18512 12640
rect 16868 12600 18512 12628
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 18598 12588 18604 12640
rect 18656 12588 18662 12640
rect 19536 12628 19564 12668
rect 20714 12628 20720 12640
rect 19536 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 21266 12628 21272 12640
rect 21223 12600 21272 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 21450 12588 21456 12640
rect 21508 12628 21514 12640
rect 21634 12628 21640 12640
rect 21508 12600 21640 12628
rect 21508 12588 21514 12600
rect 21634 12588 21640 12600
rect 21692 12628 21698 12640
rect 24765 12631 24823 12637
rect 24765 12628 24777 12631
rect 21692 12600 24777 12628
rect 21692 12588 21698 12600
rect 24765 12597 24777 12600
rect 24811 12597 24823 12631
rect 24765 12591 24823 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 4580 12396 6377 12424
rect 4580 12384 4586 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7156 12396 7481 12424
rect 7156 12384 7162 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 9858 12424 9864 12436
rect 7469 12387 7527 12393
rect 7668 12396 9864 12424
rect 4706 12356 4712 12368
rect 4448 12328 4712 12356
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 4062 12288 4068 12300
rect 1719 12260 4068 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 2130 12220 2136 12232
rect 1535 12192 2136 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2792 12229 2820 12260
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4448 12297 4476 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4203 12260 4445 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 7668 12288 7696 12396
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10594 12424 10600 12436
rect 10060 12396 10600 12424
rect 10060 12368 10088 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 11112 12396 11345 12424
rect 11112 12384 11118 12396
rect 11333 12393 11345 12396
rect 11379 12393 11391 12427
rect 11333 12387 11391 12393
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 13170 12424 13176 12436
rect 11572 12396 13176 12424
rect 11572 12384 11578 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 13872 12396 14473 12424
rect 13872 12384 13878 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 14461 12387 14519 12393
rect 14642 12384 14648 12436
rect 14700 12424 14706 12436
rect 14826 12424 14832 12436
rect 14700 12396 14832 12424
rect 14700 12384 14706 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 14918 12384 14924 12436
rect 14976 12424 14982 12436
rect 17218 12424 17224 12436
rect 14976 12396 17224 12424
rect 14976 12384 14982 12396
rect 17218 12384 17224 12396
rect 17276 12384 17282 12436
rect 17678 12384 17684 12436
rect 17736 12424 17742 12436
rect 17736 12396 18460 12424
rect 17736 12384 17742 12396
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 10042 12356 10048 12368
rect 7800 12328 10048 12356
rect 7800 12316 7806 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12356 10195 12359
rect 10778 12356 10784 12368
rect 10183 12328 10784 12356
rect 10183 12325 10195 12328
rect 10137 12319 10195 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 13630 12356 13636 12368
rect 11204 12328 13636 12356
rect 11204 12316 11210 12328
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 18432 12356 18460 12396
rect 18690 12384 18696 12436
rect 18748 12424 18754 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 18748 12396 18889 12424
rect 18748 12384 18754 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 19889 12427 19947 12433
rect 19889 12424 19901 12427
rect 19852 12396 19901 12424
rect 19852 12384 19858 12396
rect 19889 12393 19901 12396
rect 19935 12393 19947 12427
rect 20898 12424 20904 12436
rect 19889 12387 19947 12393
rect 20364 12396 20904 12424
rect 20254 12356 20260 12368
rect 14936 12328 18368 12356
rect 18432 12328 20260 12356
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 4433 12251 4491 12257
rect 4724 12260 7696 12288
rect 7944 12260 10701 12288
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 4246 12220 4252 12232
rect 2823 12192 2857 12220
rect 3160 12192 4252 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 3160 12152 3188 12192
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4724 12229 4752 12260
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5718 12180 5724 12232
rect 5776 12180 5782 12232
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 7944 12229 7972 12260
rect 10689 12257 10701 12260
rect 10735 12288 10747 12291
rect 11238 12288 11244 12300
rect 10735 12260 11244 12288
rect 10735 12257 10747 12260
rect 10689 12251 10747 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11790 12288 11796 12300
rect 11348 12260 11796 12288
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6052 12192 6837 12220
rect 6052 12180 6058 12192
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8076 12192 8800 12220
rect 8076 12180 8082 12192
rect 1964 12124 3188 12152
rect 3237 12155 3295 12161
rect 1964 12093 1992 12124
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 8202 12152 8208 12164
rect 3283 12124 8208 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 8772 12152 8800 12192
rect 8846 12180 8852 12232
rect 8904 12220 8910 12232
rect 9493 12223 9551 12229
rect 9493 12220 9505 12223
rect 8904 12192 9505 12220
rect 8904 12180 8910 12192
rect 9493 12189 9505 12192
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 11348 12220 11376 12260
rect 11790 12248 11796 12260
rect 11848 12288 11854 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11848 12260 11897 12288
rect 11848 12248 11854 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12342 12288 12348 12300
rect 12032 12260 12348 12288
rect 12032 12248 12038 12260
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 14936 12297 14964 12328
rect 13909 12291 13967 12297
rect 13909 12257 13921 12291
rect 13955 12288 13967 12291
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 13955 12260 14933 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 14752 12232 14780 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 15562 12288 15568 12300
rect 15068 12260 15568 12288
rect 15068 12248 15074 12260
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 16715 12260 18276 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 9824 12192 11376 12220
rect 9824 12180 9830 12192
rect 10704 12164 10732 12192
rect 11698 12180 11704 12232
rect 11756 12180 11762 12232
rect 12250 12220 12256 12232
rect 11808 12192 12256 12220
rect 8772 12124 9168 12152
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12084 2651 12087
rect 3786 12084 3792 12096
rect 2639 12056 3792 12084
rect 2639 12053 2651 12056
rect 2593 12047 2651 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 8018 12084 8024 12096
rect 4764 12056 8024 12084
rect 4764 12044 4770 12056
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8570 12044 8576 12096
rect 8628 12044 8634 12096
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 8812 12056 9045 12084
rect 8812 12044 8818 12056
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 9140 12084 9168 12124
rect 9674 12112 9680 12164
rect 9732 12112 9738 12164
rect 10594 12112 10600 12164
rect 10652 12112 10658 12164
rect 10686 12112 10692 12164
rect 10744 12112 10750 12164
rect 11808 12152 11836 12192
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13504 12192 14105 12220
rect 13504 12180 13510 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 15102 12220 15108 12232
rect 14875 12192 15108 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 11716 12124 11836 12152
rect 10505 12087 10563 12093
rect 10505 12084 10517 12087
rect 9140 12056 10517 12084
rect 9033 12047 9091 12053
rect 10505 12053 10517 12056
rect 10551 12084 10563 12087
rect 11716 12084 11744 12124
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12529 12155 12587 12161
rect 12529 12152 12541 12155
rect 11940 12124 12541 12152
rect 11940 12112 11946 12124
rect 12529 12121 12541 12124
rect 12575 12121 12587 12155
rect 12529 12115 12587 12121
rect 13357 12155 13415 12161
rect 13357 12121 13369 12155
rect 13403 12152 13415 12155
rect 13722 12152 13728 12164
rect 13403 12124 13728 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13722 12112 13728 12124
rect 13780 12152 13786 12164
rect 13998 12152 14004 12164
rect 13780 12124 14004 12152
rect 13780 12112 13786 12124
rect 13998 12112 14004 12124
rect 14056 12112 14062 12164
rect 14642 12112 14648 12164
rect 14700 12152 14706 12164
rect 16040 12152 16068 12183
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 18248 12229 18276 12260
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 17000 12192 17141 12220
rect 17000 12180 17006 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12189 18291 12223
rect 18340 12220 18368 12328
rect 18708 12300 18736 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 18690 12248 18696 12300
rect 18748 12248 18754 12300
rect 20364 12288 20392 12396
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 23385 12427 23443 12433
rect 23385 12424 23397 12427
rect 22796 12396 23397 12424
rect 22796 12384 22802 12396
rect 23385 12393 23397 12396
rect 23431 12393 23443 12427
rect 23385 12387 23443 12393
rect 25225 12427 25283 12433
rect 25225 12393 25237 12427
rect 25271 12424 25283 12427
rect 25314 12424 25320 12436
rect 25271 12396 25320 12424
rect 25271 12393 25283 12396
rect 25225 12387 25283 12393
rect 25314 12384 25320 12396
rect 25372 12384 25378 12436
rect 22462 12316 22468 12368
rect 22520 12356 22526 12368
rect 23474 12356 23480 12368
rect 22520 12328 23480 12356
rect 22520 12316 22526 12328
rect 23474 12316 23480 12328
rect 23532 12316 23538 12368
rect 19306 12260 20392 12288
rect 19306 12220 19334 12260
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 22646 12288 22652 12300
rect 20496 12260 22652 12288
rect 20496 12248 20502 12260
rect 22646 12248 22652 12260
rect 22704 12248 22710 12300
rect 23845 12291 23903 12297
rect 23845 12257 23857 12291
rect 23891 12288 23903 12291
rect 24210 12288 24216 12300
rect 23891 12260 24216 12288
rect 23891 12257 23903 12260
rect 23845 12251 23903 12257
rect 24210 12248 24216 12260
rect 24268 12248 24274 12300
rect 18340 12192 19334 12220
rect 18233 12183 18291 12189
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19576 12192 20085 12220
rect 19576 12180 19582 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 19978 12152 19984 12164
rect 14700 12124 15792 12152
rect 16040 12124 19984 12152
rect 14700 12112 14706 12124
rect 10551 12056 11744 12084
rect 11793 12087 11851 12093
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 11793 12053 11805 12087
rect 11839 12084 11851 12087
rect 12250 12084 12256 12096
rect 11839 12056 12256 12084
rect 11839 12053 11851 12056
rect 11793 12047 11851 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12342 12044 12348 12096
rect 12400 12084 12406 12096
rect 13446 12084 13452 12096
rect 12400 12056 13452 12084
rect 12400 12044 12406 12056
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 15010 12084 15016 12096
rect 14240 12056 15016 12084
rect 14240 12044 14246 12056
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 15764 12093 15792 12124
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 20088 12152 20116 12183
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20346 12220 20352 12232
rect 20220 12192 20352 12220
rect 20220 12180 20226 12192
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12220 24639 12223
rect 25038 12220 25044 12232
rect 24627 12192 25044 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 25038 12180 25044 12192
rect 25096 12180 25102 12232
rect 20717 12155 20775 12161
rect 20717 12152 20729 12155
rect 20088 12124 20729 12152
rect 20717 12121 20729 12124
rect 20763 12121 20775 12155
rect 22002 12152 22008 12164
rect 21942 12124 22008 12152
rect 20717 12115 20775 12121
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 15436 12056 15485 12084
rect 15436 12044 15442 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 17310 12084 17316 12096
rect 15795 12056 17316 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 17770 12044 17776 12096
rect 17828 12044 17834 12096
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 18472 12056 19349 12084
rect 18472 12044 18478 12056
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19337 12047 19395 12053
rect 19426 12044 19432 12096
rect 19484 12044 19490 12096
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 20254 12084 20260 12096
rect 19751 12056 20260 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 20254 12044 20260 12056
rect 20312 12084 20318 12096
rect 22189 12087 22247 12093
rect 22189 12084 22201 12087
rect 20312 12056 22201 12084
rect 20312 12044 20318 12056
rect 22189 12053 22201 12056
rect 22235 12053 22247 12087
rect 22189 12047 22247 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11849 1915 11883
rect 1857 11843 1915 11849
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 4798 11880 4804 11892
rect 2547 11852 4804 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 1872 11812 1900 11843
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5074 11840 5080 11892
rect 5132 11840 5138 11892
rect 9214 11880 9220 11892
rect 6104 11852 9220 11880
rect 4341 11815 4399 11821
rect 1872 11784 4292 11812
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 2038 11744 2044 11756
rect 1627 11716 2044 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2682 11704 2688 11756
rect 2740 11704 2746 11756
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3878 11744 3884 11756
rect 3375 11716 3884 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 4264 11676 4292 11784
rect 4341 11781 4353 11815
rect 4387 11812 4399 11815
rect 4433 11815 4491 11821
rect 4433 11812 4445 11815
rect 4387 11784 4445 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 4433 11781 4445 11784
rect 4479 11812 4491 11815
rect 6104 11812 6132 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 9769 11883 9827 11889
rect 9769 11880 9781 11883
rect 9640 11852 9781 11880
rect 9640 11840 9646 11852
rect 9769 11849 9781 11852
rect 9815 11849 9827 11883
rect 9769 11843 9827 11849
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 10100 11852 10149 11880
rect 10100 11840 10106 11852
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 10870 11880 10876 11892
rect 10744 11852 10876 11880
rect 10744 11840 10750 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 10965 11883 11023 11889
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11146 11880 11152 11892
rect 11011 11852 11152 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11514 11840 11520 11892
rect 11572 11840 11578 11892
rect 11793 11883 11851 11889
rect 11793 11849 11805 11883
rect 11839 11880 11851 11883
rect 11882 11880 11888 11892
rect 11839 11852 11888 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12526 11880 12532 11892
rect 12115 11852 12532 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 12676 11852 13277 11880
rect 12676 11840 12682 11852
rect 13265 11849 13277 11852
rect 13311 11849 13323 11883
rect 13265 11843 13323 11849
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13596 11852 13645 11880
rect 13596 11840 13602 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 13725 11883 13783 11889
rect 13725 11849 13737 11883
rect 13771 11880 13783 11883
rect 14274 11880 14280 11892
rect 13771 11852 14280 11880
rect 13771 11849 13783 11852
rect 13725 11843 13783 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 14550 11880 14556 11892
rect 14507 11852 14556 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 14700 11852 14933 11880
rect 14700 11840 14706 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 14921 11843 14979 11849
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 16022 11880 16028 11892
rect 15620 11852 16028 11880
rect 15620 11840 15626 11852
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 16853 11883 16911 11889
rect 16853 11849 16865 11883
rect 16899 11849 16911 11883
rect 16853 11843 16911 11849
rect 17313 11883 17371 11889
rect 17313 11849 17325 11883
rect 17359 11880 17371 11883
rect 17402 11880 17408 11892
rect 17359 11852 17408 11880
rect 17359 11849 17371 11852
rect 17313 11843 17371 11849
rect 4479 11784 6132 11812
rect 4479 11781 4491 11784
rect 4433 11775 4491 11781
rect 6638 11772 6644 11824
rect 6696 11812 6702 11824
rect 6733 11815 6791 11821
rect 6733 11812 6745 11815
rect 6696 11784 6745 11812
rect 6696 11772 6702 11784
rect 6733 11781 6745 11784
rect 6779 11781 6791 11815
rect 6733 11775 6791 11781
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 8110 11812 8116 11824
rect 6880 11784 8116 11812
rect 6880 11772 6886 11784
rect 8110 11772 8116 11784
rect 8168 11772 8174 11824
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11812 10287 11815
rect 11422 11812 11428 11824
rect 10275 11784 11428 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 11422 11772 11428 11784
rect 11480 11772 11486 11824
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 13354 11812 13360 11824
rect 11664 11784 13360 11812
rect 11664 11772 11670 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 13446 11772 13452 11824
rect 13504 11812 13510 11824
rect 16868 11812 16896 11843
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17552 11852 20760 11880
rect 17552 11840 17558 11852
rect 13504 11784 16896 11812
rect 18049 11815 18107 11821
rect 13504 11772 13510 11784
rect 18049 11781 18061 11815
rect 18095 11812 18107 11815
rect 19245 11815 19303 11821
rect 19245 11812 19257 11815
rect 18095 11784 19257 11812
rect 18095 11781 18107 11784
rect 18049 11775 18107 11781
rect 19245 11781 19257 11784
rect 19291 11812 19303 11815
rect 19426 11812 19432 11824
rect 19291 11784 19432 11812
rect 19291 11781 19303 11784
rect 19245 11775 19303 11781
rect 19426 11772 19432 11784
rect 19484 11772 19490 11824
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 20346 11812 20352 11824
rect 20220 11784 20352 11812
rect 20220 11772 20226 11784
rect 20346 11772 20352 11784
rect 20404 11772 20410 11824
rect 20732 11812 20760 11852
rect 21358 11840 21364 11892
rect 21416 11840 21422 11892
rect 21726 11812 21732 11824
rect 20732 11784 21732 11812
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 5350 11704 5356 11756
rect 5408 11704 5414 11756
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 11514 11744 11520 11756
rect 10560 11716 11520 11744
rect 10560 11704 10566 11716
rect 11514 11704 11520 11716
rect 11572 11744 11578 11756
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 11572 11716 12449 11744
rect 11572 11704 11578 11716
rect 12437 11713 12449 11716
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11744 12587 11747
rect 12618 11744 12624 11756
rect 12575 11716 12624 11744
rect 12575 11713 12587 11716
rect 12529 11707 12587 11713
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13538 11744 13544 11756
rect 13228 11716 13544 11744
rect 13228 11704 13234 11716
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13998 11704 14004 11756
rect 14056 11744 14062 11756
rect 14366 11744 14372 11756
rect 14056 11716 14372 11744
rect 14056 11704 14062 11716
rect 14366 11704 14372 11716
rect 14424 11744 14430 11756
rect 14424 11716 14780 11744
rect 14424 11704 14430 11716
rect 5902 11676 5908 11688
rect 4264 11648 5908 11676
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 5994 11636 6000 11688
rect 6052 11636 6058 11688
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 3510 11608 3516 11620
rect 2746 11580 3516 11608
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2746 11540 2774 11580
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 4522 11608 4528 11620
rect 3712 11580 4528 11608
rect 2188 11512 2774 11540
rect 3145 11543 3203 11549
rect 2188 11500 2194 11512
rect 3145 11509 3157 11543
rect 3191 11540 3203 11543
rect 3712 11540 3740 11580
rect 4522 11568 4528 11580
rect 4580 11568 4586 11620
rect 6914 11568 6920 11620
rect 6972 11568 6978 11620
rect 3191 11512 3740 11540
rect 3789 11543 3847 11549
rect 3191 11509 3203 11512
rect 3145 11503 3203 11509
rect 3789 11509 3801 11543
rect 3835 11540 3847 11543
rect 4154 11540 4160 11552
rect 3835 11512 4160 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 7098 11540 7104 11552
rect 4304 11512 7104 11540
rect 4304 11500 4310 11512
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 7392 11540 7420 11639
rect 7650 11636 7656 11688
rect 7708 11636 7714 11688
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 8662 11676 8668 11688
rect 8168 11648 8668 11676
rect 8168 11636 8174 11648
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9398 11676 9404 11688
rect 8772 11648 9404 11676
rect 8772 11552 8800 11648
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 10870 11676 10876 11688
rect 10459 11648 10876 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 12710 11636 12716 11688
rect 12768 11636 12774 11688
rect 13817 11679 13875 11685
rect 13817 11645 13829 11679
rect 13863 11645 13875 11679
rect 14182 11676 14188 11688
rect 13817 11639 13875 11645
rect 14016 11648 14188 11676
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9125 11611 9183 11617
rect 9125 11608 9137 11611
rect 8996 11580 9137 11608
rect 8996 11568 9002 11580
rect 9125 11577 9137 11580
rect 9171 11577 9183 11611
rect 9125 11571 9183 11577
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 13630 11608 13636 11620
rect 9272 11580 13636 11608
rect 9272 11568 9278 11580
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 13832 11608 13860 11639
rect 14016 11608 14044 11648
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14752 11676 14780 11716
rect 14826 11704 14832 11756
rect 14884 11704 14890 11756
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 14936 11716 15669 11744
rect 14936 11676 14964 11716
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16080 11716 17233 11744
rect 16080 11704 16086 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 18598 11744 18604 11756
rect 17221 11707 17279 11713
rect 18340 11716 18604 11744
rect 18340 11688 18368 11716
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 20254 11744 20260 11756
rect 19659 11716 20260 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 20806 11744 20812 11756
rect 20763 11716 20812 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 22097 11747 22155 11753
rect 22097 11744 22109 11747
rect 21048 11716 22109 11744
rect 21048 11704 21054 11716
rect 22097 11713 22109 11716
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 23750 11704 23756 11756
rect 23808 11744 23814 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23808 11716 23949 11744
rect 23808 11704 23814 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 14752 11648 14964 11676
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11676 17555 11679
rect 18322 11676 18328 11688
rect 17543 11648 18328 11676
rect 17543 11645 17555 11648
rect 17497 11639 17555 11645
rect 13832 11580 14044 11608
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15120 11608 15148 11639
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18564 11648 18889 11676
rect 18564 11636 18570 11648
rect 18877 11645 18889 11648
rect 18923 11676 18935 11679
rect 20622 11676 20628 11688
rect 18923 11648 20628 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 20622 11636 20628 11648
rect 20680 11636 20686 11688
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 15068 11580 15148 11608
rect 15068 11568 15074 11580
rect 8754 11540 8760 11552
rect 7392 11512 8760 11540
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 9493 11543 9551 11549
rect 9493 11509 9505 11543
rect 9539 11540 9551 11543
rect 10410 11540 10416 11552
rect 9539 11512 10416 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 16206 11540 16212 11552
rect 12032 11512 16212 11540
rect 12032 11500 12038 11512
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16298 11500 16304 11552
rect 16356 11500 16362 11552
rect 20254 11500 20260 11552
rect 20312 11500 20318 11552
rect 20346 11500 20352 11552
rect 20404 11540 20410 11552
rect 23566 11540 23572 11552
rect 20404 11512 23572 11540
rect 20404 11500 20410 11512
rect 23566 11500 23572 11512
rect 23624 11500 23630 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 3878 11336 3884 11348
rect 1627 11308 3884 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11336 4123 11339
rect 6546 11336 6552 11348
rect 4111 11308 6552 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 7469 11339 7527 11345
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 7650 11336 7656 11348
rect 7515 11308 7656 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8444 11308 8585 11336
rect 8444 11296 8450 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 9548 11308 10241 11336
rect 9548 11296 9554 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 10229 11299 10287 11305
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 11020 11308 11437 11336
rect 11020 11296 11026 11308
rect 11425 11305 11437 11308
rect 11471 11305 11483 11339
rect 11425 11299 11483 11305
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 11940 11308 13645 11336
rect 11940 11296 11946 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14366 11336 14372 11348
rect 13955 11308 14372 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14516 11308 14933 11336
rect 14516 11296 14522 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 14921 11299 14979 11305
rect 15010 11296 15016 11348
rect 15068 11336 15074 11348
rect 17494 11336 17500 11348
rect 15068 11308 17500 11336
rect 15068 11296 15074 11308
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 17862 11336 17868 11348
rect 17736 11308 17868 11336
rect 17736 11296 17742 11308
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18049 11339 18107 11345
rect 18049 11305 18061 11339
rect 18095 11336 18107 11339
rect 18966 11336 18972 11348
rect 18095 11308 18972 11336
rect 18095 11305 18107 11308
rect 18049 11299 18107 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 19334 11296 19340 11348
rect 19392 11296 19398 11348
rect 19613 11339 19671 11345
rect 19613 11305 19625 11339
rect 19659 11336 19671 11339
rect 21082 11336 21088 11348
rect 19659 11308 21088 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 22738 11296 22744 11348
rect 22796 11336 22802 11348
rect 25225 11339 25283 11345
rect 25225 11336 25237 11339
rect 22796 11308 25237 11336
rect 22796 11296 22802 11308
rect 25225 11305 25237 11308
rect 25271 11305 25283 11339
rect 25225 11299 25283 11305
rect 2593 11271 2651 11277
rect 2593 11237 2605 11271
rect 2639 11268 2651 11271
rect 4706 11268 4712 11280
rect 2639 11240 4712 11268
rect 2639 11237 2651 11240
rect 2593 11231 2651 11237
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 11606 11268 11612 11280
rect 4908 11240 11612 11268
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 2363 11172 4292 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 4062 11132 4068 11144
rect 3068 11104 4068 11132
rect 2133 11067 2191 11073
rect 2133 11033 2145 11067
rect 2179 11064 2191 11067
rect 2682 11064 2688 11076
rect 2179 11036 2688 11064
rect 2179 11033 2191 11036
rect 2133 11027 2191 11033
rect 2682 11024 2688 11036
rect 2740 11064 2746 11076
rect 3068 11064 3096 11104
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4264 11141 4292 11172
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11132 4307 11135
rect 4338 11132 4344 11144
rect 4295 11104 4344 11132
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4908 11141 4936 11240
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 11756 11240 12434 11268
rect 11756 11228 11762 11240
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 7282 11200 7288 11212
rect 5491 11172 7288 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 8202 11200 8208 11212
rect 7432 11172 8208 11200
rect 7432 11160 7438 11172
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 10318 11200 10324 11212
rect 8536 11172 10324 11200
rect 8536 11160 8542 11172
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 10870 11160 10876 11212
rect 10928 11160 10934 11212
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11790 11200 11796 11212
rect 11020 11172 11796 11200
rect 11020 11160 11026 11172
rect 11790 11160 11796 11172
rect 11848 11200 11854 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11848 11172 11989 11200
rect 11848 11160 11854 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 12406 11200 12434 11240
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 13078 11268 13084 11280
rect 12768 11240 13084 11268
rect 12768 11228 12774 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 16022 11268 16028 11280
rect 13188 11240 16028 11268
rect 13188 11200 13216 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 16114 11228 16120 11280
rect 16172 11268 16178 11280
rect 19352 11268 19380 11296
rect 16172 11240 16620 11268
rect 16172 11228 16178 11240
rect 12406 11172 13216 11200
rect 11977 11163 12035 11169
rect 13262 11160 13268 11212
rect 13320 11160 13326 11212
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 14826 11200 14832 11212
rect 13596 11172 14832 11200
rect 13596 11160 13602 11172
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 15344 11172 15393 11200
rect 15344 11160 15350 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 16206 11160 16212 11212
rect 16264 11200 16270 11212
rect 16592 11209 16620 11240
rect 17420 11240 19380 11268
rect 16577 11203 16635 11209
rect 16264 11172 16436 11200
rect 16264 11160 16270 11172
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6638 11132 6644 11144
rect 5767 11104 6644 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8386 11132 8392 11144
rect 7975 11104 8392 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 2740 11036 3096 11064
rect 3145 11067 3203 11073
rect 2740 11024 2746 11036
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 3234 11064 3240 11076
rect 3191 11036 3240 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 4798 11064 4804 11076
rect 3712 11036 4804 11064
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 2774 10996 2780 11008
rect 1912 10968 2780 10996
rect 1912 10956 1918 10968
rect 2774 10956 2780 10968
rect 2832 10996 2838 11008
rect 3712 10996 3740 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5169 11067 5227 11073
rect 5169 11064 5181 11067
rect 4908 11036 5181 11064
rect 4908 11008 4936 11036
rect 5169 11033 5181 11036
rect 5215 11033 5227 11067
rect 6840 11064 6868 11095
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8628 11104 9137 11132
rect 8628 11092 8634 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9858 11132 9864 11144
rect 9125 11095 9183 11101
rect 9232 11104 9864 11132
rect 8846 11064 8852 11076
rect 6840 11036 8852 11064
rect 5169 11027 5227 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 9232 11064 9260 11104
rect 9858 11092 9864 11104
rect 9916 11132 9922 11144
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 9916 11104 10701 11132
rect 9916 11092 9922 11104
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 13170 11132 13176 11144
rect 11931 11104 13176 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 14277 11135 14335 11141
rect 13412 11104 14228 11132
rect 13412 11092 13418 11104
rect 8996 11036 9260 11064
rect 9769 11067 9827 11073
rect 8996 11024 9002 11036
rect 9769 11033 9781 11067
rect 9815 11064 9827 11067
rect 10502 11064 10508 11076
rect 9815 11036 10508 11064
rect 9815 11033 9827 11036
rect 9769 11027 9827 11033
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11033 13047 11067
rect 12989 11027 13047 11033
rect 13081 11067 13139 11073
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 13630 11064 13636 11076
rect 13127 11036 13636 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 2832 10968 3740 10996
rect 2832 10956 2838 10968
rect 4706 10956 4712 11008
rect 4764 10956 4770 11008
rect 4890 10956 4896 11008
rect 4948 10956 4954 11008
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 6365 10999 6423 11005
rect 6365 10996 6377 10999
rect 6236 10968 6377 10996
rect 6236 10956 6242 10968
rect 6365 10965 6377 10968
rect 6411 10965 6423 10999
rect 6365 10959 6423 10965
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 10597 10999 10655 11005
rect 10597 10996 10609 10999
rect 10468 10968 10609 10996
rect 10468 10956 10474 10968
rect 10597 10965 10609 10968
rect 10643 10965 10655 10999
rect 10597 10959 10655 10965
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 11146 10996 11152 11008
rect 10744 10968 11152 10996
rect 10744 10956 10750 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 11793 10999 11851 11005
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 12158 10996 12164 11008
rect 11839 10968 12164 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12621 10999 12679 11005
rect 12621 10996 12633 10999
rect 12584 10968 12633 10996
rect 12584 10956 12590 10968
rect 12621 10965 12633 10968
rect 12667 10965 12679 10999
rect 13004 10996 13032 11027
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 14200 11064 14228 11104
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 16298 11132 16304 11144
rect 14323 11104 16304 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 16408 11141 16436 11172
rect 16577 11169 16589 11203
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 16393 11135 16451 11141
rect 16393 11101 16405 11135
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16758 11132 16764 11144
rect 16531 11104 16764 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17420 11141 17448 11240
rect 19794 11228 19800 11280
rect 19852 11268 19858 11280
rect 22189 11271 22247 11277
rect 22189 11268 22201 11271
rect 19852 11240 22201 11268
rect 19852 11228 19858 11240
rect 22189 11237 22201 11240
rect 22235 11237 22247 11271
rect 22189 11231 22247 11237
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11200 17647 11203
rect 18598 11200 18604 11212
rect 17635 11172 18604 11200
rect 17635 11169 17647 11172
rect 17589 11163 17647 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18690 11160 18696 11212
rect 18748 11160 18754 11212
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19429 11203 19487 11209
rect 19429 11200 19441 11203
rect 19024 11172 19441 11200
rect 19024 11160 19030 11172
rect 19429 11169 19441 11172
rect 19475 11169 19487 11203
rect 19429 11163 19487 11169
rect 20162 11160 20168 11212
rect 20220 11160 20226 11212
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20312 11172 24624 11200
rect 20312 11160 20318 11172
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 20809 11135 20867 11141
rect 20809 11132 20821 11135
rect 17828 11104 20821 11132
rect 17828 11092 17834 11104
rect 20809 11101 20821 11104
rect 20855 11101 20867 11135
rect 20809 11095 20867 11101
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 24596 11141 24624 11172
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 14550 11064 14556 11076
rect 13740 11036 14136 11064
rect 14200 11036 14556 11064
rect 13740 10996 13768 11036
rect 13004 10968 13768 10996
rect 14108 10996 14136 11036
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 14884 11036 15240 11064
rect 14884 11024 14890 11036
rect 15102 10996 15108 11008
rect 14108 10968 15108 10996
rect 12621 10959 12679 10965
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 15212 10996 15240 11036
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15470 11064 15476 11076
rect 15344 11036 15476 11064
rect 15344 11024 15350 11036
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 17678 11024 17684 11076
rect 17736 11064 17742 11076
rect 18417 11067 18475 11073
rect 18417 11064 18429 11067
rect 17736 11036 18429 11064
rect 17736 11024 17742 11036
rect 18417 11033 18429 11036
rect 18463 11033 18475 11067
rect 18417 11027 18475 11033
rect 18966 11024 18972 11076
rect 19024 11064 19030 11076
rect 19024 11036 20024 11064
rect 19024 11024 19030 11036
rect 16025 10999 16083 11005
rect 16025 10996 16037 10999
rect 15212 10968 16037 10996
rect 16025 10965 16037 10968
rect 16071 10965 16083 10999
rect 16025 10959 16083 10965
rect 18506 10956 18512 11008
rect 18564 10956 18570 11008
rect 19996 11005 20024 11036
rect 20346 11024 20352 11076
rect 20404 11064 20410 11076
rect 21453 11067 21511 11073
rect 21453 11064 21465 11067
rect 20404 11036 21465 11064
rect 20404 11024 20410 11036
rect 21453 11033 21465 11036
rect 21499 11033 21511 11067
rect 21453 11027 21511 11033
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 22005 11067 22063 11073
rect 22005 11064 22017 11067
rect 21692 11036 22017 11064
rect 21692 11024 21698 11036
rect 22005 11033 22017 11036
rect 22051 11033 22063 11067
rect 22005 11027 22063 11033
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 24854 11064 24860 11076
rect 23891 11036 24860 11064
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 19981 10999 20039 11005
rect 19981 10965 19993 10999
rect 20027 10965 20039 10999
rect 19981 10959 20039 10965
rect 20073 10999 20131 11005
rect 20073 10965 20085 10999
rect 20119 10996 20131 10999
rect 20162 10996 20168 11008
rect 20119 10968 20168 10996
rect 20119 10965 20131 10968
rect 20073 10959 20131 10965
rect 20162 10956 20168 10968
rect 20220 10956 20226 11008
rect 20254 10956 20260 11008
rect 20312 10996 20318 11008
rect 22278 10996 22284 11008
rect 20312 10968 22284 10996
rect 20312 10956 20318 10968
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 23658 10956 23664 11008
rect 23716 10996 23722 11008
rect 24486 10996 24492 11008
rect 23716 10968 24492 10996
rect 23716 10956 23722 10968
rect 24486 10956 24492 10968
rect 24544 10996 24550 11008
rect 25038 10996 25044 11008
rect 24544 10968 25044 10996
rect 24544 10956 24550 10968
rect 25038 10956 25044 10968
rect 25096 10956 25102 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 1854 10792 1860 10804
rect 1811 10764 1860 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 1854 10752 1860 10764
rect 1912 10752 1918 10804
rect 5258 10792 5264 10804
rect 2746 10764 5264 10792
rect 1394 10684 1400 10736
rect 1452 10724 1458 10736
rect 2746 10724 2774 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 6730 10792 6736 10804
rect 6656 10764 6736 10792
rect 1452 10696 2774 10724
rect 3421 10727 3479 10733
rect 1452 10684 1458 10696
rect 3421 10693 3433 10727
rect 3467 10724 3479 10727
rect 4706 10724 4712 10736
rect 3467 10696 4712 10724
rect 3467 10693 3479 10696
rect 3421 10687 3479 10693
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 6656 10724 6684 10764
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 8846 10752 8852 10804
rect 8904 10752 8910 10804
rect 10870 10792 10876 10804
rect 9232 10764 10876 10792
rect 4908 10696 6684 10724
rect 4908 10665 4936 10696
rect 7282 10684 7288 10736
rect 7340 10684 7346 10736
rect 7466 10684 7472 10736
rect 7524 10684 7530 10736
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 1627 10628 2881 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 2869 10625 2881 10628
rect 2915 10656 2927 10659
rect 4893 10659 4951 10665
rect 2915 10628 4016 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 2038 10548 2044 10600
rect 2096 10548 2102 10600
rect 3602 10548 3608 10600
rect 3660 10548 3666 10600
rect 2682 10412 2688 10464
rect 2740 10412 2746 10464
rect 3988 10452 4016 10628
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5902 10656 5908 10668
rect 5399 10628 5908 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 6236 10640 6684 10656
rect 6733 10643 6791 10649
rect 6733 10640 6745 10643
rect 6236 10628 6745 10640
rect 6236 10616 6242 10628
rect 6656 10612 6745 10628
rect 6733 10609 6745 10612
rect 6779 10609 6791 10643
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 8018 10656 8024 10668
rect 6972 10628 8024 10656
rect 6972 10616 6978 10628
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 9232 10656 9260 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 12713 10795 12771 10801
rect 12713 10792 12725 10795
rect 11204 10764 12725 10792
rect 11204 10752 11210 10764
rect 12713 10761 12725 10764
rect 12759 10761 12771 10795
rect 12713 10755 12771 10761
rect 13173 10795 13231 10801
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 15286 10792 15292 10804
rect 13219 10764 15292 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15804 10764 15945 10792
rect 15804 10752 15810 10764
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 9306 10684 9312 10736
rect 9364 10724 9370 10736
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 9364 10696 9597 10724
rect 9364 10684 9370 10696
rect 9585 10693 9597 10696
rect 9631 10693 9643 10727
rect 9585 10687 9643 10693
rect 10134 10684 10140 10736
rect 10192 10684 10198 10736
rect 12066 10684 12072 10736
rect 12124 10684 12130 10736
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 12176 10696 14289 10724
rect 8251 10628 9260 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 12176 10656 12204 10696
rect 14277 10693 14289 10696
rect 14323 10693 14335 10727
rect 14277 10687 14335 10693
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 15010 10724 15016 10736
rect 14424 10696 15016 10724
rect 14424 10684 14430 10696
rect 15010 10684 15016 10696
rect 15068 10724 15074 10736
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 15068 10696 15209 10724
rect 15068 10684 15074 10696
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 15948 10724 15976 10755
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 16080 10764 16681 10792
rect 16080 10752 16086 10764
rect 16669 10761 16681 10764
rect 16715 10792 16727 10795
rect 17862 10792 17868 10804
rect 16715 10764 17868 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18141 10795 18199 10801
rect 18141 10761 18153 10795
rect 18187 10792 18199 10795
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 18187 10764 21189 10792
rect 18187 10761 18199 10764
rect 18141 10755 18199 10761
rect 21177 10761 21189 10764
rect 21223 10761 21235 10795
rect 21177 10755 21235 10761
rect 21910 10752 21916 10804
rect 21968 10792 21974 10804
rect 25225 10795 25283 10801
rect 25225 10792 25237 10795
rect 21968 10764 25237 10792
rect 21968 10752 21974 10764
rect 25225 10761 25237 10764
rect 25271 10761 25283 10795
rect 25225 10755 25283 10761
rect 16206 10724 16212 10736
rect 15948 10696 16212 10724
rect 15197 10687 15255 10693
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 16482 10684 16488 10736
rect 16540 10724 16546 10736
rect 16540 10696 19472 10724
rect 16540 10684 16546 10696
rect 11112 10628 12204 10656
rect 13081 10659 13139 10665
rect 11112 10616 11118 10628
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 15470 10656 15476 10668
rect 13127 10628 15476 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 16758 10656 16764 10668
rect 16448 10628 16764 10656
rect 16448 10616 16454 10628
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17586 10656 17592 10668
rect 17083 10628 17592 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 18414 10616 18420 10668
rect 18472 10656 18478 10668
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 18472 10628 18521 10656
rect 18472 10616 18478 10628
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 19334 10656 19340 10668
rect 18509 10619 18567 10625
rect 18616 10628 19340 10656
rect 6733 10603 6791 10609
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 5994 10588 6000 10600
rect 4111 10560 6000 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 11146 10588 11152 10600
rect 9416 10560 11152 10588
rect 4709 10523 4767 10529
rect 4709 10489 4721 10523
rect 4755 10520 4767 10523
rect 4982 10520 4988 10532
rect 4755 10492 4988 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 4982 10480 4988 10492
rect 5040 10480 5046 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 9416 10520 9444 10560
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11348 10560 11928 10588
rect 6788 10492 9444 10520
rect 6788 10480 6794 10492
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 11057 10523 11115 10529
rect 11057 10520 11069 10523
rect 10928 10492 11069 10520
rect 10928 10480 10934 10492
rect 11057 10489 11069 10492
rect 11103 10520 11115 10523
rect 11348 10520 11376 10560
rect 11103 10492 11376 10520
rect 11900 10520 11928 10560
rect 13262 10548 13268 10600
rect 13320 10548 13326 10600
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13814 10588 13820 10600
rect 13412 10560 13820 10588
rect 13412 10548 13418 10560
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 14369 10591 14427 10597
rect 14369 10588 14381 10591
rect 14332 10560 14381 10588
rect 14332 10548 14338 10560
rect 14369 10557 14381 10560
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 14608 10560 15976 10588
rect 14608 10548 14614 10560
rect 13280 10520 13308 10548
rect 11900 10492 13308 10520
rect 11103 10489 11115 10492
rect 11057 10483 11115 10489
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 13596 10492 15577 10520
rect 13596 10480 13602 10492
rect 15565 10489 15577 10492
rect 15611 10489 15623 10523
rect 15948 10520 15976 10560
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 16132 10520 16160 10551
rect 17310 10548 17316 10600
rect 17368 10588 17374 10600
rect 18616 10597 18644 10628
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 17368 10560 18613 10588
rect 17368 10548 17374 10560
rect 18601 10557 18613 10560
rect 18647 10557 18659 10591
rect 18601 10551 18659 10557
rect 18785 10591 18843 10597
rect 18785 10557 18797 10591
rect 18831 10588 18843 10591
rect 19150 10588 19156 10600
rect 18831 10560 19156 10588
rect 18831 10557 18843 10560
rect 18785 10551 18843 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 16482 10520 16488 10532
rect 15948 10492 16488 10520
rect 15565 10483 15623 10489
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 18506 10520 18512 10532
rect 17604 10492 18512 10520
rect 5074 10452 5080 10464
rect 3988 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 5776 10424 6009 10452
rect 5776 10412 5782 10424
rect 5997 10421 6009 10424
rect 6043 10421 6055 10455
rect 5997 10415 6055 10421
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6914 10452 6920 10464
rect 6595 10424 6920 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 7926 10452 7932 10464
rect 7800 10424 7932 10452
rect 7800 10412 7806 10424
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 10226 10452 10232 10464
rect 8076 10424 10232 10452
rect 8076 10412 8082 10424
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 10376 10424 11713 10452
rect 10376 10412 10382 10424
rect 11701 10421 11713 10424
rect 11747 10452 11759 10455
rect 11790 10452 11796 10464
rect 11747 10424 11796 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11940 10424 12173 10452
rect 11940 10412 11946 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13814 10452 13820 10464
rect 13228 10424 13820 10452
rect 13228 10412 13234 10424
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 13906 10412 13912 10464
rect 13964 10412 13970 10464
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 14826 10452 14832 10464
rect 14332 10424 14832 10452
rect 14332 10412 14338 10424
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 14918 10412 14924 10464
rect 14976 10452 14982 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14976 10424 15025 10452
rect 14976 10412 14982 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 17604 10452 17632 10492
rect 18506 10480 18512 10492
rect 18564 10520 18570 10532
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 18564 10492 19257 10520
rect 18564 10480 18570 10492
rect 19245 10489 19257 10492
rect 19291 10489 19303 10523
rect 19245 10483 19303 10489
rect 15160 10424 17632 10452
rect 15160 10412 15166 10424
rect 17678 10412 17684 10464
rect 17736 10412 17742 10464
rect 19444 10452 19472 10696
rect 20254 10684 20260 10736
rect 20312 10684 20318 10736
rect 22370 10684 22376 10736
rect 22428 10684 22434 10736
rect 23290 10684 23296 10736
rect 23348 10684 23354 10736
rect 25038 10684 25044 10736
rect 25096 10684 25102 10736
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 20346 10656 20352 10668
rect 19659 10628 20352 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10656 22155 10659
rect 22554 10656 22560 10668
rect 22143 10628 22560 10656
rect 22143 10625 22155 10628
rect 22097 10619 22155 10625
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22704 10628 23029 10656
rect 22704 10616 22710 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23017 10619 23075 10625
rect 24394 10616 24400 10668
rect 24452 10616 24458 10668
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10557 21327 10591
rect 21269 10551 21327 10557
rect 19702 10480 19708 10532
rect 19760 10520 19766 10532
rect 21284 10520 21312 10551
rect 22278 10548 22284 10600
rect 22336 10588 22342 10600
rect 25409 10591 25467 10597
rect 25409 10588 25421 10591
rect 22336 10560 25421 10588
rect 22336 10548 22342 10560
rect 25409 10557 25421 10560
rect 25455 10557 25467 10591
rect 25409 10551 25467 10557
rect 22370 10520 22376 10532
rect 19760 10492 22376 10520
rect 19760 10480 19766 10492
rect 22370 10480 22376 10492
rect 22428 10480 22434 10532
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 19444 10424 20729 10452
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 20717 10415 20775 10421
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 24765 10455 24823 10461
rect 24765 10452 24777 10455
rect 23532 10424 24777 10452
rect 23532 10412 23538 10424
rect 24765 10421 24777 10424
rect 24811 10421 24823 10455
rect 24765 10415 24823 10421
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 2961 10251 3019 10257
rect 2961 10217 2973 10251
rect 3007 10248 3019 10251
rect 5902 10248 5908 10260
rect 3007 10220 5908 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6052 10220 7880 10248
rect 6052 10208 6058 10220
rect 1581 10183 1639 10189
rect 1581 10149 1593 10183
rect 1627 10149 1639 10183
rect 1581 10143 1639 10149
rect 2225 10183 2283 10189
rect 2225 10149 2237 10183
rect 2271 10180 2283 10183
rect 3973 10183 4031 10189
rect 2271 10152 3924 10180
rect 2271 10149 2283 10152
rect 2225 10143 2283 10149
rect 1394 10072 1400 10124
rect 1452 10072 1458 10124
rect 1596 10112 1624 10143
rect 3896 10112 3924 10152
rect 3973 10149 3985 10183
rect 4019 10180 4031 10183
rect 4246 10180 4252 10192
rect 4019 10152 4252 10180
rect 4019 10149 4031 10152
rect 3973 10143 4031 10149
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 7742 10180 7748 10192
rect 4632 10152 7748 10180
rect 4632 10112 4660 10152
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 7852 10180 7880 10220
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8444 10220 8585 10248
rect 8444 10208 8450 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 9122 10248 9128 10260
rect 8720 10220 9128 10248
rect 8720 10208 8726 10220
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9232 10220 10640 10248
rect 9232 10180 9260 10220
rect 7852 10152 9260 10180
rect 1596 10084 3832 10112
rect 3896 10084 4660 10112
rect 4709 10115 4767 10121
rect 1412 10044 1440 10072
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 1412 10016 1777 10044
rect 1765 10013 1777 10016
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 3418 10044 3424 10056
rect 2455 10016 3424 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 1394 9936 1400 9988
rect 1452 9976 1458 9988
rect 2424 9976 2452 10007
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 1452 9948 2452 9976
rect 2777 9979 2835 9985
rect 1452 9936 1458 9948
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 3234 9976 3240 9988
rect 2823 9948 3240 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 3804 9908 3832 10084
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 4755 10084 6377 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 8478 10112 8484 10124
rect 6365 10075 6423 10081
rect 6472 10084 8484 10112
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4172 9976 4200 10007
rect 5718 10004 5724 10056
rect 5776 10004 5782 10056
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 6472 10044 6500 10084
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 9398 10112 9404 10124
rect 9171 10084 9404 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9398 10072 9404 10084
rect 9456 10112 9462 10124
rect 9766 10112 9772 10124
rect 9456 10084 9772 10112
rect 9456 10072 9462 10084
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 5960 10016 6500 10044
rect 6825 10047 6883 10053
rect 5960 10004 5966 10016
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 7282 10044 7288 10056
rect 6871 10016 7288 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 9030 10044 9036 10056
rect 7975 10016 9036 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 10612 10044 10640 10220
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 11241 10251 11299 10257
rect 11241 10248 11253 10251
rect 10744 10220 11253 10248
rect 10744 10208 10750 10220
rect 11241 10217 11253 10220
rect 11287 10217 11299 10251
rect 11241 10211 11299 10217
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11572 10220 11805 10248
rect 11572 10208 11578 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 12216 10220 13001 10248
rect 12216 10208 12222 10220
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 14274 10248 14280 10260
rect 12989 10211 13047 10217
rect 13096 10220 14280 10248
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 11204 10152 11437 10180
rect 11204 10140 11210 10152
rect 11425 10149 11437 10152
rect 11471 10180 11483 10183
rect 12526 10180 12532 10192
rect 11471 10152 12532 10180
rect 11471 10149 11483 10152
rect 11425 10143 11483 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 13096 10180 13124 10220
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 14724 10251 14782 10257
rect 14724 10217 14736 10251
rect 14770 10248 14782 10251
rect 14770 10220 15792 10248
rect 14770 10217 14782 10220
rect 14724 10211 14782 10217
rect 14182 10180 14188 10192
rect 12768 10152 13124 10180
rect 13464 10152 14188 10180
rect 12768 10140 12774 10152
rect 10870 10072 10876 10124
rect 10928 10072 10934 10124
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 11514 10112 11520 10124
rect 11296 10084 11520 10112
rect 11296 10072 11302 10084
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 11664 10084 12357 10112
rect 11664 10072 11670 10084
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 10612 10016 12173 10044
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 13464 10044 13492 10152
rect 14182 10140 14188 10152
rect 14240 10180 14246 10192
rect 14366 10180 14372 10192
rect 14240 10152 14372 10180
rect 14240 10140 14246 10152
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 15764 10180 15792 10220
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 15896 10220 16681 10248
rect 15896 10208 15902 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17184 10220 17785 10248
rect 17184 10208 17190 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 19702 10248 19708 10260
rect 17920 10220 19708 10248
rect 17920 10208 17926 10220
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 20036 10220 20085 10248
rect 20036 10208 20042 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 20073 10211 20131 10217
rect 20714 10208 20720 10260
rect 20772 10208 20778 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 22833 10251 22891 10257
rect 22833 10248 22845 10251
rect 20956 10220 22845 10248
rect 20956 10208 20962 10220
rect 22833 10217 22845 10220
rect 22879 10217 22891 10251
rect 22833 10211 22891 10217
rect 25225 10251 25283 10257
rect 25225 10217 25237 10251
rect 25271 10248 25283 10251
rect 25682 10248 25688 10260
rect 25271 10220 25688 10248
rect 25271 10217 25283 10220
rect 25225 10211 25283 10217
rect 25682 10208 25688 10220
rect 25740 10208 25746 10260
rect 16850 10180 16856 10192
rect 15764 10152 16856 10180
rect 16850 10140 16856 10152
rect 16908 10140 16914 10192
rect 18690 10140 18696 10192
rect 18748 10180 18754 10192
rect 20732 10180 20760 10208
rect 18748 10152 20760 10180
rect 18748 10140 18754 10152
rect 22370 10140 22376 10192
rect 22428 10140 22434 10192
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 13648 10084 17172 10112
rect 13403 10016 13492 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 4172 9948 7052 9976
rect 4982 9908 4988 9920
rect 3804 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 5442 9908 5448 9920
rect 5307 9880 5448 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 7024 9908 7052 9948
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 7156 9948 9413 9976
rect 7156 9936 7162 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 9401 9939 9459 9945
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9548 9948 9812 9976
rect 9548 9936 9554 9948
rect 7190 9908 7196 9920
rect 7024 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 9582 9908 9588 9920
rect 7515 9880 9588 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9784 9908 9812 9948
rect 10134 9936 10140 9988
rect 10192 9936 10198 9988
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 10836 9948 12265 9976
rect 10836 9936 10842 9948
rect 12253 9945 12265 9948
rect 12299 9945 12311 9979
rect 12253 9939 12311 9945
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 13648 9976 13676 10084
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 13872 10016 14473 10044
rect 13872 10004 13878 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15870 10016 16589 10044
rect 14461 10007 14519 10013
rect 16577 10013 16589 10016
rect 16623 10044 16635 10047
rect 16758 10044 16764 10056
rect 16623 10016 16764 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17144 10053 17172 10084
rect 19242 10072 19248 10124
rect 19300 10112 19306 10124
rect 23474 10112 23480 10124
rect 19300 10084 23480 10112
rect 19300 10072 19306 10084
rect 23474 10072 23480 10084
rect 23532 10072 23538 10124
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17678 10004 17684 10056
rect 17736 10044 17742 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 17736 10016 18245 10044
rect 17736 10004 17742 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19429 10047 19487 10053
rect 19429 10044 19441 10047
rect 18380 10016 19441 10044
rect 18380 10004 18386 10016
rect 19429 10013 19441 10016
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 20622 10004 20628 10056
rect 20680 10004 20686 10056
rect 22002 10004 22008 10056
rect 22060 10004 22066 10056
rect 23198 10004 23204 10056
rect 23256 10004 23262 10056
rect 24302 10004 24308 10056
rect 24360 10044 24366 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24360 10016 24593 10044
rect 24360 10004 24366 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 14734 9976 14740 9988
rect 13596 9948 13676 9976
rect 14108 9948 14740 9976
rect 13596 9936 13602 9948
rect 11054 9908 11060 9920
rect 9784 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 11572 9880 13461 9908
rect 11572 9868 11578 9880
rect 13449 9877 13461 9880
rect 13495 9908 13507 9911
rect 14108 9908 14136 9948
rect 14734 9936 14740 9948
rect 14792 9936 14798 9988
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 20901 9979 20959 9985
rect 20901 9976 20913 9979
rect 16448 9948 20913 9976
rect 16448 9936 16454 9948
rect 20901 9945 20913 9948
rect 20947 9945 20959 9979
rect 20901 9939 20959 9945
rect 13495 9880 14136 9908
rect 14185 9911 14243 9917
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 14185 9877 14197 9911
rect 14231 9908 14243 9911
rect 14550 9908 14556 9920
rect 14231 9880 14556 9908
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 14550 9868 14556 9880
rect 14608 9908 14614 9920
rect 14826 9908 14832 9920
rect 14608 9880 14832 9908
rect 14608 9868 14614 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16114 9908 16120 9920
rect 15712 9880 16120 9908
rect 15712 9868 15718 9880
rect 16114 9868 16120 9880
rect 16172 9908 16178 9920
rect 16209 9911 16267 9917
rect 16209 9908 16221 9911
rect 16172 9880 16221 9908
rect 16172 9868 16178 9880
rect 16209 9877 16221 9880
rect 16255 9877 16267 9911
rect 16209 9871 16267 9877
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 17862 9908 17868 9920
rect 16816 9880 17868 9908
rect 16816 9868 16822 9880
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18322 9868 18328 9920
rect 18380 9908 18386 9920
rect 18690 9908 18696 9920
rect 18380 9880 18696 9908
rect 18380 9868 18386 9880
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 18877 9911 18935 9917
rect 18877 9877 18889 9911
rect 18923 9908 18935 9911
rect 18966 9908 18972 9920
rect 18923 9880 18972 9908
rect 18923 9877 18935 9880
rect 18877 9871 18935 9877
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 22278 9908 22284 9920
rect 19484 9880 22284 9908
rect 19484 9868 19490 9880
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 22830 9868 22836 9920
rect 22888 9908 22894 9920
rect 23293 9911 23351 9917
rect 23293 9908 23305 9911
rect 22888 9880 23305 9908
rect 22888 9868 22894 9880
rect 23293 9877 23305 9880
rect 23339 9877 23351 9911
rect 23293 9871 23351 9877
rect 23842 9868 23848 9920
rect 23900 9868 23906 9920
rect 24026 9868 24032 9920
rect 24084 9868 24090 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 4080 9676 4844 9704
rect 1397 9639 1455 9645
rect 1397 9605 1409 9639
rect 1443 9636 1455 9639
rect 1443 9608 2820 9636
rect 1443 9605 1455 9608
rect 1397 9599 1455 9605
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 1544 9540 2145 9568
rect 1544 9528 1550 9540
rect 2133 9537 2145 9540
rect 2179 9568 2191 9571
rect 2222 9568 2228 9580
rect 2179 9540 2228 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2792 9577 2820 9608
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 4080 9636 4108 9676
rect 3344 9608 4108 9636
rect 4157 9639 4215 9645
rect 2785 9571 2843 9577
rect 2785 9537 2797 9571
rect 2831 9568 2843 9571
rect 3344 9568 3372 9608
rect 4157 9605 4169 9639
rect 4203 9636 4215 9639
rect 4430 9636 4436 9648
rect 4203 9608 4436 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4580 9608 4721 9636
rect 4580 9596 4586 9608
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 4816 9636 4844 9676
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 8202 9704 8208 9716
rect 5316 9676 8208 9704
rect 5316 9664 5322 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9030 9664 9036 9716
rect 9088 9704 9094 9716
rect 10870 9704 10876 9716
rect 9088 9676 10876 9704
rect 9088 9664 9094 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 12158 9704 12164 9716
rect 11296 9676 12164 9704
rect 11296 9664 11302 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 13449 9707 13507 9713
rect 12308 9676 13308 9704
rect 12308 9664 12314 9676
rect 6178 9636 6184 9648
rect 4816 9608 6184 9636
rect 4709 9599 4767 9605
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 7282 9596 7288 9648
rect 7340 9596 7346 9648
rect 7650 9596 7656 9648
rect 7708 9636 7714 9648
rect 9398 9636 9404 9648
rect 7708 9608 9404 9636
rect 7708 9596 7714 9608
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 11333 9639 11391 9645
rect 2831 9540 3372 9568
rect 3973 9571 4031 9577
rect 2831 9537 2843 9540
rect 2785 9531 2843 9537
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 1854 9500 1860 9512
rect 1719 9472 1860 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 3988 9500 4016 9531
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4304 9540 5365 9568
rect 4304 9528 4310 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9568 6055 9571
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6043 9540 6653 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 10336 9568 10364 9622
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 12434 9636 12440 9648
rect 11379 9608 12440 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13280 9636 13308 9676
rect 13449 9673 13461 9707
rect 13495 9704 13507 9707
rect 13998 9704 14004 9716
rect 13495 9676 14004 9704
rect 13495 9673 13507 9676
rect 13449 9667 13507 9673
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 14553 9707 14611 9713
rect 14553 9673 14565 9707
rect 14599 9673 14611 9707
rect 14553 9667 14611 9673
rect 16868 9676 17080 9704
rect 14568 9636 14596 9667
rect 13280 9608 14596 9636
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 14700 9608 15056 9636
rect 14700 9596 14706 9608
rect 10410 9568 10416 9580
rect 10336 9540 10416 9568
rect 7745 9531 7803 9537
rect 7558 9500 7564 9512
rect 3988 9472 7564 9500
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 1949 9435 2007 9441
rect 1949 9432 1961 9435
rect 1360 9404 1961 9432
rect 1360 9392 1366 9404
rect 1949 9401 1961 9404
rect 1995 9401 2007 9435
rect 1949 9395 2007 9401
rect 2314 9392 2320 9444
rect 2372 9432 2378 9444
rect 7374 9432 7380 9444
rect 2372 9404 7380 9432
rect 2372 9392 2378 9404
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 7760 9432 7788 9531
rect 10410 9528 10416 9540
rect 10468 9568 10474 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10468 9540 10885 9568
rect 10468 9528 10474 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 13504 9540 14044 9568
rect 13504 9528 13510 9540
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8812 9472 8861 9500
rect 8812 9460 8818 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 9824 9472 11713 9500
rect 9824 9460 9830 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12618 9500 12624 9512
rect 12023 9472 12624 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 7760 9404 8984 9432
rect 2590 9324 2596 9376
rect 2648 9324 2654 9376
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4522 9364 4528 9376
rect 4120 9336 4528 9364
rect 4120 9324 4126 9336
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 4982 9364 4988 9376
rect 4847 9336 4988 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 7708 9336 8401 9364
rect 7708 9324 7714 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8956 9364 8984 9404
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10410 9432 10416 9444
rect 10192 9404 10416 9432
rect 10192 9392 10198 9404
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 11606 9432 11612 9444
rect 10612 9404 11612 9432
rect 10612 9373 10640 9404
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 8956 9336 10609 9364
rect 8389 9327 8447 9333
rect 10597 9333 10609 9336
rect 10643 9333 10655 9367
rect 10597 9327 10655 9333
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11514 9364 11520 9376
rect 11195 9336 11520 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11716 9364 11744 9463
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13228 9472 13921 9500
rect 13228 9460 13234 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 14016 9500 14044 9540
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14424 9540 14933 9568
rect 14424 9528 14430 9540
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 15028 9568 15056 9608
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 15896 9608 16129 9636
rect 15896 9596 15902 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 16206 9596 16212 9648
rect 16264 9636 16270 9648
rect 16868 9636 16896 9676
rect 16264 9608 16896 9636
rect 16264 9596 16270 9608
rect 16942 9596 16948 9648
rect 17000 9596 17006 9648
rect 17052 9636 17080 9676
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 20530 9704 20536 9716
rect 17276 9676 20536 9704
rect 17276 9664 17282 9676
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 24026 9704 24032 9716
rect 20772 9676 24032 9704
rect 20772 9664 20778 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 18414 9636 18420 9648
rect 17052 9608 18420 9636
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 19613 9639 19671 9645
rect 19613 9605 19625 9639
rect 19659 9636 19671 9639
rect 19886 9636 19892 9648
rect 19659 9608 19892 9636
rect 19659 9605 19671 9608
rect 19613 9599 19671 9605
rect 19886 9596 19892 9608
rect 19944 9596 19950 9648
rect 19978 9596 19984 9648
rect 20036 9636 20042 9648
rect 20036 9608 23980 9636
rect 20036 9596 20042 9608
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 15028 9540 18153 9568
rect 14921 9531 14979 9537
rect 18141 9537 18153 9540
rect 18187 9568 18199 9571
rect 18187 9540 18460 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 14016 9472 14780 9500
rect 13909 9463 13967 9469
rect 14752 9444 14780 9472
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14884 9472 15025 9500
rect 14884 9460 14890 9472
rect 15013 9469 15025 9472
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 15102 9460 15108 9512
rect 15160 9460 15166 9512
rect 15212 9472 17540 9500
rect 13722 9432 13728 9444
rect 13372 9404 13728 9432
rect 12710 9364 12716 9376
rect 11716 9336 12716 9364
rect 12710 9324 12716 9336
rect 12768 9364 12774 9376
rect 13372 9364 13400 9404
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14182 9432 14188 9444
rect 14056 9404 14188 9432
rect 14056 9392 14062 9404
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 15120 9432 15148 9460
rect 14792 9404 15148 9432
rect 14792 9392 14798 9404
rect 12768 9336 13400 9364
rect 12768 9324 12774 9336
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 15212 9364 15240 9472
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9432 15715 9435
rect 16114 9432 16120 9444
rect 15703 9404 16120 9432
rect 15703 9401 15715 9404
rect 15657 9395 15715 9401
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 16298 9392 16304 9444
rect 16356 9392 16362 9444
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 16816 9404 17417 9432
rect 16816 9392 16822 9404
rect 17405 9401 17417 9404
rect 17451 9401 17463 9435
rect 17512 9432 17540 9472
rect 17586 9460 17592 9512
rect 17644 9500 17650 9512
rect 18230 9500 18236 9512
rect 17644 9472 18236 9500
rect 17644 9460 17650 9472
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18322 9460 18328 9512
rect 18380 9460 18386 9512
rect 18432 9500 18460 9540
rect 18966 9528 18972 9580
rect 19024 9528 19030 9580
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9568 20315 9571
rect 20346 9568 20352 9580
rect 20303 9540 20352 9568
rect 20303 9537 20315 9540
rect 20257 9531 20315 9537
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 20456 9540 22109 9568
rect 19610 9500 19616 9512
rect 18432 9472 19616 9500
rect 19610 9460 19616 9472
rect 19668 9460 19674 9512
rect 20456 9432 20484 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23658 9568 23664 9580
rect 22796 9540 23664 9568
rect 22796 9528 22802 9540
rect 23658 9528 23664 9540
rect 23716 9528 23722 9580
rect 23952 9577 23980 9608
rect 23937 9571 23995 9577
rect 23937 9537 23949 9571
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 22278 9500 22284 9512
rect 21315 9472 22284 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 23290 9460 23296 9512
rect 23348 9460 23354 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 17512 9404 20484 9432
rect 17405 9395 17463 9401
rect 20990 9392 20996 9444
rect 21048 9432 21054 9444
rect 21542 9432 21548 9444
rect 21048 9404 21548 9432
rect 21048 9392 21054 9404
rect 21542 9392 21548 9404
rect 21600 9392 21606 9444
rect 13504 9336 15240 9364
rect 13504 9324 13510 9336
rect 17034 9324 17040 9376
rect 17092 9324 17098 9376
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 17494 9364 17500 9376
rect 17184 9336 17500 9364
rect 17184 9324 17190 9336
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17770 9324 17776 9376
rect 17828 9324 17834 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 22462 9364 22468 9376
rect 19024 9336 22468 9364
rect 19024 9324 19030 9336
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 2501 9163 2559 9169
rect 2501 9129 2513 9163
rect 2547 9160 2559 9163
rect 4706 9160 4712 9172
rect 2547 9132 4712 9160
rect 2547 9129 2559 9132
rect 2501 9123 2559 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 8938 9160 8944 9172
rect 6696 9132 8944 9160
rect 6696 9120 6702 9132
rect 8938 9120 8944 9132
rect 8996 9160 9002 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8996 9132 9045 9160
rect 8996 9120 9002 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 9180 9132 11161 9160
rect 9180 9120 9186 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 12066 9160 12072 9172
rect 11747 9132 12072 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 12618 9120 12624 9172
rect 12676 9120 12682 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 14737 9163 14795 9169
rect 14737 9160 14749 9163
rect 13688 9132 14749 9160
rect 13688 9120 13694 9132
rect 14737 9129 14749 9132
rect 14783 9129 14795 9163
rect 14737 9123 14795 9129
rect 15930 9120 15936 9172
rect 15988 9120 15994 9172
rect 19337 9163 19395 9169
rect 19337 9160 19349 9163
rect 16408 9132 19349 9160
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 3510 9092 3516 9104
rect 1903 9064 3516 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 6362 9092 6368 9104
rect 4120 9064 6368 9092
rect 4120 9052 4126 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 11790 9092 11796 9104
rect 10284 9064 11796 9092
rect 10284 9052 10290 9064
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 16022 9092 16028 9104
rect 12860 9064 16028 9092
rect 12860 9052 12866 9064
rect 16022 9052 16028 9064
rect 16080 9052 16086 9104
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 7469 9027 7527 9033
rect 2464 8996 7328 9024
rect 2464 8984 2470 8996
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2038 8956 2044 8968
rect 1728 8928 2044 8956
rect 1728 8916 1734 8928
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2682 8916 2688 8968
rect 2740 8916 2746 8968
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 4614 8916 4620 8968
rect 4672 8916 4678 8968
rect 5258 8916 5264 8968
rect 5316 8916 5322 8968
rect 5718 8916 5724 8968
rect 5776 8916 5782 8968
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 7190 8956 7196 8968
rect 6871 8928 7196 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 3237 8891 3295 8897
rect 3237 8888 3249 8891
rect 1636 8860 3249 8888
rect 1636 8848 1642 8860
rect 3237 8857 3249 8860
rect 3283 8857 3295 8891
rect 6730 8888 6736 8900
rect 3237 8851 3295 8857
rect 3896 8860 6736 8888
rect 1486 8780 1492 8832
rect 1544 8780 1550 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3896 8820 3924 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7300 8888 7328 8996
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 8846 9024 8852 9036
rect 7515 8996 8852 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 10594 9024 10600 9036
rect 9416 8996 10600 9024
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8294 8956 8300 8968
rect 7975 8928 8300 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9416 8965 9444 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 12342 9024 12348 9036
rect 11204 8996 12348 9024
rect 11204 8984 11210 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 13814 9024 13820 9036
rect 12584 8996 13820 9024
rect 12584 8984 12590 8996
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 14056 8996 14105 9024
rect 14056 8984 14062 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 14240 8996 14381 9024
rect 14240 8984 14246 8996
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 14918 9024 14924 9036
rect 14516 8996 14924 9024
rect 14516 8984 14522 8996
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 9024 15439 9027
rect 15562 9024 15568 9036
rect 15427 8996 15568 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9548 8928 10437 8956
rect 9548 8916 9554 8928
rect 10226 8888 10232 8900
rect 7300 8860 10232 8888
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 10409 8888 10437 8928
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12434 8956 12440 8968
rect 12023 8928 12440 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8956 13139 8959
rect 16114 8956 16120 8968
rect 13127 8928 16120 8956
rect 13127 8925 13139 8928
rect 13081 8919 13139 8925
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 11238 8888 11244 8900
rect 10409 8860 11244 8888
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 12308 8860 14136 8888
rect 12308 8848 12314 8860
rect 3200 8792 3924 8820
rect 3200 8780 3206 8792
rect 3970 8780 3976 8832
rect 4028 8780 4034 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 6365 8823 6423 8829
rect 6365 8820 6377 8823
rect 5408 8792 6377 8820
rect 5408 8780 5414 8792
rect 6365 8789 6377 8792
rect 6411 8789 6423 8823
rect 6365 8783 6423 8789
rect 8570 8780 8576 8832
rect 8628 8780 8634 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10045 8823 10103 8829
rect 10045 8820 10057 8823
rect 9732 8792 10057 8820
rect 9732 8780 9738 8792
rect 10045 8789 10057 8792
rect 10091 8789 10103 8823
rect 10045 8783 10103 8789
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 10836 8792 11437 8820
rect 10836 8780 10842 8792
rect 11425 8789 11437 8792
rect 11471 8820 11483 8823
rect 13630 8820 13636 8832
rect 11471 8792 13636 8820
rect 11471 8789 11483 8792
rect 11425 8783 11483 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13722 8780 13728 8832
rect 13780 8780 13786 8832
rect 14108 8820 14136 8860
rect 14182 8848 14188 8900
rect 14240 8888 14246 8900
rect 16408 8897 16436 9132
rect 19337 9129 19349 9132
rect 19383 9160 19395 9163
rect 19794 9160 19800 9172
rect 19383 9132 19800 9160
rect 19383 9129 19395 9132
rect 19337 9123 19395 9129
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 21637 9163 21695 9169
rect 21637 9160 21649 9163
rect 19904 9132 21649 9160
rect 19150 9052 19156 9104
rect 19208 9092 19214 9104
rect 19904 9092 19932 9132
rect 21637 9129 21649 9132
rect 21683 9129 21695 9163
rect 21637 9123 21695 9129
rect 25222 9120 25228 9172
rect 25280 9120 25286 9172
rect 19208 9064 19932 9092
rect 19208 9052 19214 9064
rect 16482 8984 16488 9036
rect 16540 8984 16546 9036
rect 17402 8984 17408 9036
rect 17460 8984 17466 9036
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 19889 9027 19947 9033
rect 19889 9024 19901 9027
rect 17552 8996 19901 9024
rect 17552 8984 17558 8996
rect 19889 8993 19901 8996
rect 19935 9024 19947 9027
rect 20622 9024 20628 9036
rect 19935 8996 20628 9024
rect 19935 8993 19947 8996
rect 19889 8987 19947 8993
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 22281 9027 22339 9033
rect 22281 8993 22293 9027
rect 22327 9024 22339 9027
rect 22646 9024 22652 9036
rect 22327 8996 22652 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 17126 8916 17132 8968
rect 17184 8916 17190 8968
rect 21910 8956 21916 8968
rect 21298 8928 21916 8956
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22002 8916 22008 8968
rect 22060 8956 22066 8968
rect 22296 8956 22324 8987
rect 22646 8984 22652 8996
rect 22704 8984 22710 9036
rect 22060 8928 22324 8956
rect 24581 8959 24639 8965
rect 22060 8916 22066 8928
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 24670 8956 24676 8968
rect 24627 8928 24676 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 16393 8891 16451 8897
rect 16393 8888 16405 8891
rect 14240 8860 16405 8888
rect 14240 8848 14246 8860
rect 16393 8857 16405 8860
rect 16439 8857 16451 8891
rect 16393 8851 16451 8857
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 17494 8888 17500 8900
rect 16540 8860 17500 8888
rect 16540 8848 16546 8860
rect 15102 8820 15108 8832
rect 14108 8792 15108 8820
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 16206 8820 16212 8832
rect 15252 8792 16212 8820
rect 15252 8780 15258 8792
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16301 8823 16359 8829
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 16592 8820 16620 8860
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 17954 8848 17960 8900
rect 18012 8848 18018 8900
rect 18690 8848 18696 8900
rect 18748 8888 18754 8900
rect 20165 8891 20223 8897
rect 20165 8888 20177 8891
rect 18748 8860 20177 8888
rect 18748 8848 18754 8860
rect 20165 8857 20177 8860
rect 20211 8857 20223 8891
rect 21928 8888 21956 8916
rect 21928 8860 22048 8888
rect 20165 8851 20223 8857
rect 16347 8792 16620 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 18877 8823 18935 8829
rect 18877 8820 18889 8823
rect 16724 8792 18889 8820
rect 16724 8780 16730 8792
rect 18877 8789 18889 8792
rect 18923 8789 18935 8823
rect 18877 8783 18935 8789
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 19429 8823 19487 8829
rect 19429 8820 19441 8823
rect 19300 8792 19441 8820
rect 19300 8780 19306 8792
rect 19429 8789 19441 8792
rect 19475 8789 19487 8823
rect 19429 8783 19487 8789
rect 19610 8780 19616 8832
rect 19668 8820 19674 8832
rect 21913 8823 21971 8829
rect 21913 8820 21925 8823
rect 19668 8792 21925 8820
rect 19668 8780 19674 8792
rect 21913 8789 21925 8792
rect 21959 8789 21971 8823
rect 22020 8820 22048 8860
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 22557 8891 22615 8897
rect 22557 8888 22569 8891
rect 22152 8860 22569 8888
rect 22152 8848 22158 8860
rect 22557 8857 22569 8860
rect 22603 8857 22615 8891
rect 22557 8851 22615 8857
rect 22756 8860 23046 8888
rect 22756 8832 22784 8860
rect 22738 8820 22744 8832
rect 22020 8792 22744 8820
rect 21913 8783 21971 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 22830 8780 22836 8832
rect 22888 8820 22894 8832
rect 24029 8823 24087 8829
rect 24029 8820 24041 8823
rect 22888 8792 24041 8820
rect 22888 8780 22894 8792
rect 24029 8789 24041 8792
rect 24075 8789 24087 8823
rect 24029 8783 24087 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 3142 8616 3148 8628
rect 1811 8588 3148 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3329 8619 3387 8625
rect 3329 8585 3341 8619
rect 3375 8616 3387 8619
rect 6822 8616 6828 8628
rect 3375 8588 6828 8616
rect 3375 8585 3387 8588
rect 3329 8579 3387 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7190 8576 7196 8628
rect 7248 8576 7254 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7742 8616 7748 8628
rect 7524 8588 7748 8616
rect 7524 8576 7530 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8294 8576 8300 8628
rect 8352 8576 8358 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 8404 8588 10977 8616
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 1535 8520 2728 8548
rect 1535 8517 1547 8520
rect 1489 8511 1547 8517
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1946 8480 1952 8492
rect 1636 8452 1952 8480
rect 1636 8440 1642 8452
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2700 8480 2728 8520
rect 2774 8508 2780 8560
rect 2832 8548 2838 8560
rect 3237 8551 3295 8557
rect 3237 8548 3249 8551
rect 2832 8520 3249 8548
rect 2832 8508 2838 8520
rect 3237 8517 3249 8520
rect 3283 8517 3295 8551
rect 3237 8511 3295 8517
rect 3786 8508 3792 8560
rect 3844 8548 3850 8560
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3844 8520 3985 8548
rect 3844 8508 3850 8520
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 3973 8511 4031 8517
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 4709 8551 4767 8557
rect 4709 8548 4721 8551
rect 4212 8520 4721 8548
rect 4212 8508 4218 8520
rect 4709 8517 4721 8520
rect 4755 8517 4767 8551
rect 4709 8511 4767 8517
rect 4893 8551 4951 8557
rect 4893 8517 4905 8551
rect 4939 8548 4951 8551
rect 5902 8548 5908 8560
rect 4939 8520 5908 8548
rect 4939 8517 4951 8520
rect 4893 8511 4951 8517
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 6362 8508 6368 8560
rect 6420 8548 6426 8560
rect 6638 8548 6644 8560
rect 6420 8520 6644 8548
rect 6420 8508 6426 8520
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 7558 8508 7564 8560
rect 7616 8548 7622 8560
rect 8404 8548 8432 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 12434 8576 12440 8628
rect 12492 8576 12498 8628
rect 13814 8616 13820 8628
rect 13556 8588 13820 8616
rect 7616 8520 8432 8548
rect 7616 8508 7622 8520
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 8628 8520 9045 8548
rect 8628 8508 8634 8520
rect 9033 8517 9045 8520
rect 9079 8517 9091 8551
rect 13556 8548 13584 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 13964 8588 14013 8616
rect 13964 8576 13970 8588
rect 14001 8585 14013 8588
rect 14047 8585 14059 8619
rect 14001 8579 14059 8585
rect 14366 8576 14372 8628
rect 14424 8576 14430 8628
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 16758 8616 16764 8628
rect 15160 8588 16764 8616
rect 15160 8576 15166 8588
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8616 17279 8619
rect 18322 8616 18328 8628
rect 17267 8588 18328 8616
rect 17267 8585 17279 8588
rect 17221 8579 17279 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 20438 8576 20444 8628
rect 20496 8616 20502 8628
rect 20496 8588 23980 8616
rect 20496 8576 20502 8588
rect 9033 8511 9091 8517
rect 10336 8520 13584 8548
rect 4062 8480 4068 8492
rect 2700 8452 4068 8480
rect 2501 8443 2559 8449
rect 2516 8412 2544 8443
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 6549 8483 6607 8489
rect 6196 8452 6500 8480
rect 4157 8415 4215 8421
rect 2516 8384 4108 8412
rect 2682 8304 2688 8356
rect 2740 8304 2746 8356
rect 4080 8344 4108 8384
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 6196 8412 6224 8452
rect 4203 8384 6224 8412
rect 6472 8412 6500 8452
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 7466 8480 7472 8492
rect 6595 8452 7472 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 8386 8412 8392 8424
rect 6472 8384 8392 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8754 8372 8760 8424
rect 8812 8372 8818 8424
rect 10336 8412 10364 8520
rect 13630 8508 13636 8560
rect 13688 8548 13694 8560
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 13688 8520 14473 8548
rect 13688 8508 13694 8520
rect 14461 8517 14473 8520
rect 14507 8548 14519 8551
rect 14642 8548 14648 8560
rect 14507 8520 14648 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 15562 8508 15568 8560
rect 15620 8548 15626 8560
rect 16206 8548 16212 8560
rect 15620 8520 16212 8548
rect 15620 8508 15626 8520
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 16942 8508 16948 8560
rect 17000 8548 17006 8560
rect 17402 8548 17408 8560
rect 17000 8520 17408 8548
rect 17000 8508 17006 8520
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 17494 8508 17500 8560
rect 17552 8548 17558 8560
rect 19242 8548 19248 8560
rect 17552 8520 19248 8548
rect 17552 8508 17558 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 19429 8551 19487 8557
rect 19429 8517 19441 8551
rect 19475 8548 19487 8551
rect 21542 8548 21548 8560
rect 19475 8520 21548 8548
rect 19475 8517 19487 8520
rect 19429 8511 19487 8517
rect 21542 8508 21548 8520
rect 21600 8508 21606 8560
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 8864 8384 10364 8412
rect 5350 8344 5356 8356
rect 4080 8316 5356 8344
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5718 8344 5724 8356
rect 5552 8316 5724 8344
rect 1118 8236 1124 8288
rect 1176 8276 1182 8288
rect 3878 8276 3884 8288
rect 1176 8248 3884 8276
rect 1176 8236 1182 8248
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5552 8276 5580 8316
rect 5718 8304 5724 8316
rect 5776 8344 5782 8356
rect 5776 8316 6132 8344
rect 5776 8304 5782 8316
rect 5316 8248 5580 8276
rect 5316 8236 5322 8248
rect 5994 8236 6000 8288
rect 6052 8236 6058 8288
rect 6104 8276 6132 8316
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 8864 8344 8892 8384
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 11808 8412 11836 8443
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12492 8452 12909 8480
rect 12492 8440 12498 8452
rect 12897 8449 12909 8452
rect 12943 8480 12955 8483
rect 12943 8452 14320 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 10744 8384 11836 8412
rect 10744 8372 10750 8384
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13630 8412 13636 8424
rect 13320 8384 13636 8412
rect 13320 8372 13326 8384
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13872 8384 13921 8412
rect 13872 8372 13878 8384
rect 13909 8381 13921 8384
rect 13955 8412 13967 8415
rect 14292 8412 14320 8452
rect 14476 8452 15700 8480
rect 14476 8412 14504 8452
rect 13955 8384 14228 8412
rect 14292 8384 14504 8412
rect 14553 8415 14611 8421
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 7432 8316 8892 8344
rect 10505 8347 10563 8353
rect 7432 8304 7438 8316
rect 10505 8313 10517 8347
rect 10551 8344 10563 8347
rect 10594 8344 10600 8356
rect 10551 8316 10600 8344
rect 10551 8313 10563 8316
rect 10505 8307 10563 8313
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 10928 8316 12204 8344
rect 10928 8304 10934 8316
rect 9214 8276 9220 8288
rect 6104 8248 9220 8276
rect 9214 8236 9220 8248
rect 9272 8276 9278 8288
rect 12066 8276 12072 8288
rect 9272 8248 12072 8276
rect 9272 8236 9278 8248
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12176 8276 12204 8316
rect 12802 8304 12808 8356
rect 12860 8344 12866 8356
rect 13446 8344 13452 8356
rect 12860 8316 13452 8344
rect 12860 8304 12866 8316
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 13538 8304 13544 8356
rect 13596 8304 13602 8356
rect 14200 8344 14228 8384
rect 14553 8381 14565 8415
rect 14599 8381 14611 8415
rect 14553 8375 14611 8381
rect 14366 8344 14372 8356
rect 13740 8316 13952 8344
rect 14200 8316 14372 8344
rect 13740 8276 13768 8316
rect 13924 8288 13952 8316
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 14458 8304 14464 8356
rect 14516 8344 14522 8356
rect 14568 8344 14596 8375
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 15194 8412 15200 8424
rect 14700 8384 15200 8412
rect 14700 8372 14706 8384
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 14734 8344 14740 8356
rect 14516 8316 14740 8344
rect 14516 8304 14522 8316
rect 14734 8304 14740 8316
rect 14792 8304 14798 8356
rect 14826 8304 14832 8356
rect 14884 8344 14890 8356
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 14884 8316 15025 8344
rect 14884 8304 14890 8316
rect 15013 8313 15025 8316
rect 15059 8313 15071 8347
rect 15013 8307 15071 8313
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 15528 8316 15577 8344
rect 15528 8304 15534 8316
rect 15565 8313 15577 8316
rect 15611 8313 15623 8347
rect 15672 8344 15700 8452
rect 15930 8440 15936 8492
rect 15988 8440 15994 8492
rect 17957 8483 18015 8489
rect 17957 8480 17969 8483
rect 16040 8452 17969 8480
rect 15746 8372 15752 8424
rect 15804 8412 15810 8424
rect 16040 8421 16068 8452
rect 17957 8449 17969 8452
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15804 8384 16037 8412
rect 15804 8372 15810 8384
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 16206 8372 16212 8424
rect 16264 8372 16270 8424
rect 17218 8372 17224 8424
rect 17276 8412 17282 8424
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 17276 8384 17325 8412
rect 17276 8372 17282 8384
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 16666 8344 16672 8356
rect 15672 8316 16672 8344
rect 15565 8307 15623 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 17678 8344 17684 8356
rect 16899 8316 17684 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 17972 8344 18000 8443
rect 18432 8412 18460 8443
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 18748 8452 20085 8480
rect 18748 8440 18754 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 23952 8489 23980 8588
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 22097 8483 22155 8489
rect 22097 8480 22109 8483
rect 20220 8452 22109 8480
rect 20220 8440 20226 8452
rect 22097 8449 22109 8452
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 18966 8412 18972 8424
rect 18432 8384 18972 8412
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 21174 8412 21180 8424
rect 19300 8384 21180 8412
rect 19300 8372 19306 8384
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 22370 8412 22376 8424
rect 21315 8384 22376 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 22370 8372 22376 8384
rect 22428 8372 22434 8424
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 24854 8412 24860 8424
rect 23339 8384 24860 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 20254 8344 20260 8356
rect 17972 8316 20260 8344
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 12176 8248 13768 8276
rect 13906 8236 13912 8288
rect 13964 8236 13970 8288
rect 18782 8236 18788 8288
rect 18840 8276 18846 8288
rect 18966 8276 18972 8288
rect 18840 8248 18972 8276
rect 18840 8236 18846 8248
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 20438 8276 20444 8288
rect 19392 8248 20444 8276
rect 19392 8236 19398 8248
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2406 8072 2412 8084
rect 1912 8044 2412 8072
rect 1912 8032 1918 8044
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 4982 8072 4988 8084
rect 4847 8044 4988 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5258 8032 5264 8084
rect 5316 8032 5322 8084
rect 5442 8032 5448 8084
rect 5500 8032 5506 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 7098 8072 7104 8084
rect 6411 8044 7104 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7466 8032 7472 8084
rect 7524 8032 7530 8084
rect 9030 8072 9036 8084
rect 7852 8044 9036 8072
rect 1210 7964 1216 8016
rect 1268 8004 1274 8016
rect 1578 8004 1584 8016
rect 1268 7976 1584 8004
rect 1268 7964 1274 7976
rect 1578 7964 1584 7976
rect 1636 7964 1642 8016
rect 3421 8007 3479 8013
rect 3421 7973 3433 8007
rect 3467 8004 3479 8007
rect 3510 8004 3516 8016
rect 3467 7976 3516 8004
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 3510 7964 3516 7976
rect 3568 7964 3574 8016
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7936 1547 7939
rect 3142 7936 3148 7948
rect 1535 7908 3148 7936
rect 1535 7905 1547 7908
rect 1489 7899 1547 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 7852 7936 7880 8044
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 10134 8072 10140 8084
rect 9180 8044 10140 8072
rect 9180 8032 9186 8044
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 11698 8072 11704 8084
rect 11195 8044 11704 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 19610 8072 19616 8084
rect 12124 8044 19616 8072
rect 12124 8032 12130 8044
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 20438 8032 20444 8084
rect 20496 8032 20502 8084
rect 25225 8075 25283 8081
rect 25225 8041 25237 8075
rect 25271 8072 25283 8075
rect 25590 8072 25596 8084
rect 25271 8044 25596 8072
rect 25271 8041 25283 8044
rect 25225 8035 25283 8041
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 12250 8004 12256 8016
rect 7984 7976 9812 8004
rect 7984 7964 7990 7976
rect 9674 7936 9680 7948
rect 3252 7908 7880 7936
rect 7944 7908 9680 7936
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 3252 7877 3280 7908
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 2464 7840 2513 7868
rect 2464 7828 2470 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 4614 7868 4620 7880
rect 3237 7831 3295 7837
rect 3804 7840 4620 7868
rect 2685 7803 2743 7809
rect 2685 7769 2697 7803
rect 2731 7800 2743 7803
rect 3804 7800 3832 7840
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4706 7828 4712 7880
rect 4764 7828 4770 7880
rect 7944 7877 7972 7908
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 2731 7772 3832 7800
rect 2731 7769 2743 7772
rect 2685 7763 2743 7769
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 1765 7735 1823 7741
rect 1765 7732 1777 7735
rect 1728 7704 1777 7732
rect 1728 7692 1734 7704
rect 1765 7701 1777 7704
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 3973 7735 4031 7741
rect 3973 7701 3985 7735
rect 4019 7732 4031 7735
rect 4706 7732 4712 7744
rect 4019 7704 4712 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 5736 7732 5764 7831
rect 6840 7800 6868 7831
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8352 7840 9045 7868
rect 8352 7828 8358 7840
rect 9033 7837 9045 7840
rect 9079 7868 9091 7871
rect 9122 7868 9128 7880
rect 9079 7840 9128 7868
rect 9079 7837 9091 7840
rect 9033 7831 9091 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9364 7840 9413 7868
rect 9364 7828 9370 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 9784 7800 9812 7976
rect 10060 7976 12256 8004
rect 10060 7877 10088 7976
rect 12250 7964 12256 7976
rect 12308 8004 12314 8016
rect 12308 7976 14872 8004
rect 12308 7964 12314 7976
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11296 7908 11621 7936
rect 11296 7896 11302 7908
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7936 11851 7939
rect 12434 7936 12440 7948
rect 11839 7908 12440 7936
rect 11839 7905 11851 7908
rect 11793 7899 11851 7905
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 12894 7896 12900 7948
rect 12952 7896 12958 7948
rect 13446 7896 13452 7948
rect 13504 7936 13510 7948
rect 14642 7936 14648 7948
rect 13504 7908 14648 7936
rect 13504 7896 13510 7908
rect 14642 7896 14648 7908
rect 14700 7896 14706 7948
rect 14844 7945 14872 7976
rect 15286 7964 15292 8016
rect 15344 8004 15350 8016
rect 15657 8007 15715 8013
rect 15657 8004 15669 8007
rect 15344 7976 15669 8004
rect 15344 7964 15350 7976
rect 15657 7973 15669 7976
rect 15703 7973 15715 8007
rect 15657 7967 15715 7973
rect 16758 7964 16764 8016
rect 16816 8004 16822 8016
rect 16853 8007 16911 8013
rect 16853 8004 16865 8007
rect 16816 7976 16865 8004
rect 16816 7964 16822 7976
rect 16853 7973 16865 7976
rect 16899 7973 16911 8007
rect 19334 8004 19340 8016
rect 16853 7967 16911 7973
rect 16960 7976 19340 8004
rect 14829 7939 14887 7945
rect 14829 7905 14841 7939
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15381 7939 15439 7945
rect 15381 7936 15393 7939
rect 14976 7908 15393 7936
rect 14976 7896 14982 7908
rect 15381 7905 15393 7908
rect 15427 7905 15439 7939
rect 15381 7899 15439 7905
rect 16206 7896 16212 7948
rect 16264 7896 16270 7948
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 16960 7936 16988 7976
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 19429 8007 19487 8013
rect 19429 7973 19441 8007
rect 19475 8004 19487 8007
rect 24026 8004 24032 8016
rect 19475 7976 24032 8004
rect 19475 7973 19487 7976
rect 19429 7967 19487 7973
rect 24026 7964 24032 7976
rect 24084 7964 24090 8016
rect 19886 7936 19892 7948
rect 16448 7908 16988 7936
rect 17052 7908 19892 7936
rect 16448 7896 16454 7908
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10192 7840 11652 7868
rect 10192 7828 10198 7840
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 6840 7772 9352 7800
rect 9784 7772 11529 7800
rect 8478 7732 8484 7744
rect 5736 7704 8484 7732
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 8846 7732 8852 7744
rect 8619 7704 8852 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 9324 7732 9352 7772
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 11624 7800 11652 7840
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 12216 7840 13737 7868
rect 12216 7828 12222 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 17052 7877 17080 7908
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20073 7939 20131 7945
rect 20073 7905 20085 7939
rect 20119 7936 20131 7939
rect 20254 7936 20260 7948
rect 20119 7908 20260 7936
rect 20119 7905 20131 7908
rect 20073 7899 20131 7905
rect 20254 7896 20260 7908
rect 20312 7936 20318 7948
rect 22830 7936 22836 7948
rect 20312 7908 22836 7936
rect 20312 7896 20318 7908
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24854 7936 24860 7948
rect 23891 7908 24860 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 13964 7840 16037 7868
rect 13964 7828 13970 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17494 7828 17500 7880
rect 17552 7828 17558 7880
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 17644 7840 20821 7868
rect 17644 7828 17650 7840
rect 20809 7837 20821 7840
rect 20855 7837 20867 7871
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 20809 7831 20867 7837
rect 20916 7840 22661 7868
rect 11624 7772 13676 7800
rect 11517 7763 11575 7769
rect 10962 7732 10968 7744
rect 9324 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 12345 7735 12403 7741
rect 12345 7732 12357 7735
rect 11848 7704 12357 7732
rect 11848 7692 11854 7704
rect 12345 7701 12357 7704
rect 12391 7701 12403 7735
rect 12345 7695 12403 7701
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 12584 7704 12725 7732
rect 12584 7692 12590 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 12713 7695 12771 7701
rect 12802 7692 12808 7744
rect 12860 7692 12866 7744
rect 13538 7692 13544 7744
rect 13596 7692 13602 7744
rect 13648 7732 13676 7772
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14737 7803 14795 7809
rect 14737 7800 14749 7803
rect 13872 7772 14749 7800
rect 13872 7760 13878 7772
rect 14737 7769 14749 7772
rect 14783 7769 14795 7803
rect 14737 7763 14795 7769
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 15160 7772 16129 7800
rect 15160 7760 15166 7772
rect 16117 7769 16129 7772
rect 16163 7800 16175 7803
rect 17402 7800 17408 7812
rect 16163 7772 17408 7800
rect 16163 7769 16175 7772
rect 16117 7763 16175 7769
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 18693 7803 18751 7809
rect 18693 7769 18705 7803
rect 18739 7800 18751 7803
rect 19058 7800 19064 7812
rect 18739 7772 19064 7800
rect 18739 7769 18751 7772
rect 18693 7763 18751 7769
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 19610 7800 19616 7812
rect 19168 7772 19616 7800
rect 14182 7732 14188 7744
rect 13648 7704 14188 7732
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14274 7692 14280 7744
rect 14332 7692 14338 7744
rect 14642 7692 14648 7744
rect 14700 7692 14706 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 19168 7732 19196 7772
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 19794 7760 19800 7812
rect 19852 7760 19858 7812
rect 19978 7760 19984 7812
rect 20036 7800 20042 7812
rect 20916 7800 20944 7840
rect 22649 7837 22661 7840
rect 22695 7837 22707 7871
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 22649 7831 22707 7837
rect 24412 7840 24593 7868
rect 20036 7772 20944 7800
rect 22005 7803 22063 7809
rect 20036 7760 20042 7772
rect 22005 7769 22017 7803
rect 22051 7800 22063 7803
rect 22462 7800 22468 7812
rect 22051 7772 22468 7800
rect 22051 7769 22063 7772
rect 22005 7763 22063 7769
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 24412 7744 24440 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 16632 7704 19196 7732
rect 16632 7692 16638 7704
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19702 7732 19708 7744
rect 19392 7704 19708 7732
rect 19392 7692 19398 7704
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 19886 7692 19892 7744
rect 19944 7692 19950 7744
rect 24394 7692 24400 7744
rect 24452 7692 24458 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 1820 7500 2329 7528
rect 1820 7488 1826 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 5258 7528 5264 7540
rect 2648 7500 5264 7528
rect 2648 7488 2654 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6822 7528 6828 7540
rect 6043 7500 6828 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 10318 7528 10324 7540
rect 6932 7500 10324 7528
rect 3418 7420 3424 7472
rect 3476 7460 3482 7472
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 3476 7432 3709 7460
rect 3476 7420 3482 7432
rect 3697 7429 3709 7432
rect 3743 7429 3755 7463
rect 3697 7423 3755 7429
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 5718 7460 5724 7472
rect 3936 7432 5724 7460
rect 3936 7420 3942 7432
rect 5718 7420 5724 7432
rect 5776 7420 5782 7472
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2682 7392 2688 7404
rect 1719 7364 2688 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2774 7352 2780 7404
rect 2832 7352 2838 7404
rect 3970 7392 3976 7404
rect 2884 7364 3976 7392
rect 2884 7324 2912 7364
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4120 7364 4261 7392
rect 4120 7352 4126 7364
rect 4249 7361 4261 7364
rect 4295 7392 4307 7395
rect 4338 7392 4344 7404
rect 4295 7364 4344 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 5994 7392 6000 7404
rect 5399 7364 6000 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6932 7401 6960 7500
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 10410 7488 10416 7540
rect 10468 7528 10474 7540
rect 10468 7500 10732 7528
rect 10468 7488 10474 7500
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 8665 7463 8723 7469
rect 8665 7460 8677 7463
rect 8628 7432 8677 7460
rect 8628 7420 8634 7432
rect 8665 7429 8677 7432
rect 8711 7460 8723 7463
rect 9490 7460 9496 7472
rect 8711 7432 9496 7460
rect 8711 7429 8723 7432
rect 8665 7423 8723 7429
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 10704 7460 10732 7500
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 12618 7528 12624 7540
rect 11020 7500 12624 7528
rect 11020 7488 11026 7500
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13372 7500 18184 7528
rect 10626 7432 11284 7460
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 11256 7401 11284 7432
rect 12360 7432 12848 7460
rect 12360 7404 12388 7432
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7524 7364 8033 7392
rect 7524 7352 7530 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11287 7364 11621 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 11609 7361 11621 7364
rect 11655 7392 11667 7395
rect 11793 7395 11851 7401
rect 11793 7392 11805 7395
rect 11655 7364 11805 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 11793 7361 11805 7364
rect 11839 7392 11851 7395
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11839 7364 11989 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11977 7361 11989 7364
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12342 7352 12348 7404
rect 12400 7352 12406 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 12492 7364 12633 7392
rect 12492 7352 12498 7364
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 2746 7296 2912 7324
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 2746 7256 2774 7296
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 7006 7324 7012 7336
rect 3200 7296 7012 7324
rect 3200 7284 3206 7296
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8812 7296 9137 7324
rect 8812 7284 8818 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 10134 7324 10140 7336
rect 9447 7296 10140 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 2372 7228 2774 7256
rect 2372 7216 2378 7228
rect 2866 7216 2872 7268
rect 2924 7256 2930 7268
rect 3510 7256 3516 7268
rect 2924 7228 3516 7256
rect 2924 7216 2930 7228
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 3970 7216 3976 7268
rect 4028 7256 4034 7268
rect 4982 7256 4988 7268
rect 4028 7228 4988 7256
rect 4028 7216 4034 7228
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 5040 7228 6040 7256
rect 5040 7216 5046 7228
rect 6012 7200 6040 7228
rect 3418 7148 3424 7200
rect 3476 7148 3482 7200
rect 4890 7148 4896 7200
rect 4948 7148 4954 7200
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 6052 7160 6377 7188
rect 6052 7148 6058 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6638 7148 6644 7200
rect 6696 7148 6702 7200
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 9140 7188 9168 7287
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 12820 7333 12848 7432
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 11388 7296 12725 7324
rect 11388 7284 11394 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 10410 7216 10416 7268
rect 10468 7256 10474 7268
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 10468 7228 10885 7256
rect 10468 7216 10474 7228
rect 10873 7225 10885 7228
rect 10919 7256 10931 7259
rect 12894 7256 12900 7268
rect 10919 7228 12900 7256
rect 10919 7225 10931 7228
rect 10873 7219 10931 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 9398 7188 9404 7200
rect 9140 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11790 7188 11796 7200
rect 11480 7160 11796 7188
rect 11480 7148 11486 7160
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12253 7191 12311 7197
rect 12253 7188 12265 7191
rect 12032 7160 12265 7188
rect 12032 7148 12038 7160
rect 12253 7157 12265 7160
rect 12299 7157 12311 7191
rect 12253 7151 12311 7157
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 13372 7188 13400 7500
rect 15562 7460 15568 7472
rect 14950 7432 15568 7460
rect 15562 7420 15568 7432
rect 15620 7420 15626 7472
rect 16206 7420 16212 7472
rect 16264 7460 16270 7472
rect 16301 7463 16359 7469
rect 16301 7460 16313 7463
rect 16264 7432 16313 7460
rect 16264 7420 16270 7432
rect 16301 7429 16313 7432
rect 16347 7429 16359 7463
rect 17313 7463 17371 7469
rect 17313 7460 17325 7463
rect 16301 7423 16359 7429
rect 16408 7432 17325 7460
rect 15654 7352 15660 7404
rect 15712 7352 15718 7404
rect 15930 7352 15936 7404
rect 15988 7392 15994 7404
rect 16408 7392 16436 7432
rect 17313 7429 17325 7432
rect 17359 7429 17371 7463
rect 17313 7423 17371 7429
rect 17402 7420 17408 7472
rect 17460 7460 17466 7472
rect 18156 7469 18184 7500
rect 18524 7500 19288 7528
rect 17497 7463 17555 7469
rect 17497 7460 17509 7463
rect 17460 7432 17509 7460
rect 17460 7420 17466 7432
rect 17497 7429 17509 7432
rect 17543 7429 17555 7463
rect 17497 7423 17555 7429
rect 18141 7463 18199 7469
rect 18141 7429 18153 7463
rect 18187 7429 18199 7463
rect 18141 7423 18199 7429
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 18524 7460 18552 7500
rect 18288 7432 18630 7460
rect 18288 7420 18294 7432
rect 19260 7404 19288 7500
rect 22066 7500 23612 7528
rect 22066 7460 22094 7500
rect 19444 7432 22094 7460
rect 15988 7364 16436 7392
rect 15988 7352 15994 7364
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16816 7364 17049 7392
rect 16816 7352 16822 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 13449 7327 13507 7333
rect 13449 7293 13461 7327
rect 13495 7293 13507 7327
rect 13449 7287 13507 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 17402 7324 17408 7336
rect 13771 7296 17408 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 12400 7160 13400 7188
rect 13464 7188 13492 7287
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 16022 7256 16028 7268
rect 14752 7228 16028 7256
rect 14752 7188 14780 7228
rect 16022 7216 16028 7228
rect 16080 7256 16086 7268
rect 17126 7256 17132 7268
rect 16080 7228 17132 7256
rect 16080 7216 16086 7228
rect 17126 7216 17132 7228
rect 17184 7256 17190 7268
rect 17880 7256 17908 7287
rect 18598 7284 18604 7336
rect 18656 7324 18662 7336
rect 18874 7324 18880 7336
rect 18656 7296 18880 7324
rect 18656 7284 18662 7296
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 17184 7228 17908 7256
rect 17184 7216 17190 7228
rect 13464 7160 14780 7188
rect 12400 7148 12406 7160
rect 15194 7148 15200 7200
rect 15252 7148 15258 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16390 7188 16396 7200
rect 16264 7160 16396 7188
rect 16264 7148 16270 7160
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 16853 7191 16911 7197
rect 16853 7188 16865 7191
rect 16632 7160 16865 7188
rect 16632 7148 16638 7160
rect 16853 7157 16865 7160
rect 16899 7157 16911 7191
rect 16853 7151 16911 7157
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 19444 7188 19472 7432
rect 22738 7420 22744 7472
rect 22796 7420 22802 7472
rect 23584 7460 23612 7500
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 24029 7531 24087 7537
rect 24029 7528 24041 7531
rect 23992 7500 24041 7528
rect 23992 7488 23998 7500
rect 24029 7497 24041 7500
rect 24075 7497 24087 7531
rect 24029 7491 24087 7497
rect 24213 7463 24271 7469
rect 24213 7460 24225 7463
rect 23584 7432 24225 7460
rect 24213 7429 24225 7432
rect 24259 7460 24271 7463
rect 24259 7432 24440 7460
rect 24259 7429 24271 7432
rect 24213 7423 24271 7429
rect 19610 7352 19616 7404
rect 19668 7392 19674 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 19668 7364 20085 7392
rect 19668 7352 19674 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 24412 7401 24440 7432
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 22646 7324 22652 7336
rect 21315 7296 22652 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 22646 7284 22652 7296
rect 22704 7284 22710 7336
rect 24118 7284 24124 7336
rect 24176 7324 24182 7336
rect 24673 7327 24731 7333
rect 24673 7324 24685 7327
rect 24176 7296 24685 7324
rect 24176 7284 24182 7296
rect 24673 7293 24685 7296
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 23753 7259 23811 7265
rect 23753 7225 23765 7259
rect 23799 7256 23811 7259
rect 23842 7256 23848 7268
rect 23799 7228 23848 7256
rect 23799 7225 23811 7228
rect 23753 7219 23811 7225
rect 23842 7216 23848 7228
rect 23900 7256 23906 7268
rect 25314 7256 25320 7268
rect 23900 7228 25320 7256
rect 23900 7216 23906 7228
rect 25314 7216 25320 7228
rect 25372 7216 25378 7268
rect 17920 7160 19472 7188
rect 17920 7148 17926 7160
rect 19610 7148 19616 7200
rect 19668 7148 19674 7200
rect 22094 7148 22100 7200
rect 22152 7188 22158 7200
rect 22262 7191 22320 7197
rect 22262 7188 22274 7191
rect 22152 7160 22274 7188
rect 22152 7148 22158 7160
rect 22262 7157 22274 7160
rect 22308 7157 22320 7191
rect 22262 7151 22320 7157
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 4614 6944 4620 6996
rect 4672 6984 4678 6996
rect 8938 6984 8944 6996
rect 4672 6956 8944 6984
rect 4672 6944 4678 6956
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 10870 6984 10876 6996
rect 10704 6956 10876 6984
rect 2130 6876 2136 6928
rect 2188 6916 2194 6928
rect 2866 6916 2872 6928
rect 2188 6888 2872 6916
rect 2188 6876 2194 6888
rect 2866 6876 2872 6888
rect 2924 6876 2930 6928
rect 5074 6876 5080 6928
rect 5132 6916 5138 6928
rect 5132 6888 5764 6916
rect 5132 6876 5138 6888
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 2314 6848 2320 6860
rect 1627 6820 2320 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 5626 6848 5632 6860
rect 2884 6820 5632 6848
rect 1118 6740 1124 6792
rect 1176 6780 1182 6792
rect 2884 6789 2912 6820
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5736 6848 5764 6888
rect 6546 6876 6552 6928
rect 6604 6916 6610 6928
rect 10704 6916 10732 6956
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 12342 6984 12348 6996
rect 11112 6956 12348 6984
rect 11112 6944 11118 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 19610 6984 19616 6996
rect 12676 6956 19616 6984
rect 12676 6944 12682 6956
rect 19610 6944 19616 6956
rect 19668 6944 19674 6996
rect 16758 6916 16764 6928
rect 6604 6888 10732 6916
rect 12728 6888 16764 6916
rect 6604 6876 6610 6888
rect 5736 6820 6592 6848
rect 6564 6792 6592 6820
rect 9214 6808 9220 6860
rect 9272 6808 9278 6860
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 9456 6820 10609 6848
rect 9456 6808 9462 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 12308 6820 12357 6848
rect 12308 6808 12314 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 12728 6857 12756 6888
rect 16758 6876 16764 6888
rect 16816 6876 16822 6928
rect 17494 6876 17500 6928
rect 17552 6916 17558 6928
rect 19794 6916 19800 6928
rect 17552 6888 19800 6916
rect 17552 6876 17558 6888
rect 19794 6876 19800 6888
rect 19852 6876 19858 6928
rect 19886 6876 19892 6928
rect 19944 6916 19950 6928
rect 19944 6888 20024 6916
rect 19944 6876 19950 6888
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12676 6820 12725 6848
rect 12676 6808 12682 6820
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 13998 6848 14004 6860
rect 12713 6811 12771 6817
rect 13004 6820 14004 6848
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1176 6752 1961 6780
rect 1176 6740 1182 6752
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 1949 6743 2007 6749
rect 2056 6752 2605 6780
rect 566 6672 572 6724
rect 624 6712 630 6724
rect 1302 6712 1308 6724
rect 624 6684 1308 6712
rect 624 6672 630 6684
rect 1302 6672 1308 6684
rect 1360 6712 1366 6724
rect 2056 6712 2084 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 5537 6783 5595 6789
rect 4120 6752 5120 6780
rect 4120 6740 4126 6752
rect 1360 6684 2084 6712
rect 2133 6715 2191 6721
rect 1360 6672 1366 6684
rect 2133 6681 2145 6715
rect 2179 6712 2191 6715
rect 4982 6712 4988 6724
rect 2179 6684 4988 6712
rect 2179 6681 2191 6684
rect 2133 6675 2191 6681
rect 4982 6672 4988 6684
rect 5040 6672 5046 6724
rect 5092 6712 5120 6752
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5583 6752 5733 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 5721 6749 5733 6752
rect 5767 6780 5779 6783
rect 5902 6780 5908 6792
rect 5767 6752 5908 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8754 6780 8760 6792
rect 7975 6752 8760 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 6270 6712 6276 6724
rect 5092 6684 6276 6712
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 6840 6712 6868 6743
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 8904 6752 9505 6780
rect 8904 6740 8910 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 11974 6740 11980 6792
rect 12032 6740 12038 6792
rect 13004 6780 13032 6820
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6848 15715 6851
rect 15746 6848 15752 6860
rect 15703 6820 15752 6848
rect 15703 6817 15715 6820
rect 15657 6811 15715 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 18506 6848 18512 6860
rect 15988 6820 18512 6848
rect 15988 6808 15994 6820
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 18598 6808 18604 6860
rect 18656 6808 18662 6860
rect 19996 6857 20024 6888
rect 19981 6851 20039 6857
rect 19981 6817 19993 6851
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 20128 6820 20453 6848
rect 20128 6808 20134 6820
rect 20441 6817 20453 6820
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 25317 6851 25375 6857
rect 25317 6817 25329 6851
rect 25363 6848 25375 6851
rect 25498 6848 25504 6860
rect 25363 6820 25504 6848
rect 25363 6817 25375 6820
rect 25317 6811 25375 6817
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 12176 6752 13032 6780
rect 13081 6783 13139 6789
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 6840 6684 8585 6712
rect 8573 6681 8585 6684
rect 8619 6681 8631 6715
rect 10778 6712 10784 6724
rect 8573 6675 8631 6681
rect 9232 6684 10784 6712
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4120 6616 4629 6644
rect 4120 6604 4126 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 5077 6647 5135 6653
rect 5077 6613 5089 6647
rect 5123 6644 5135 6647
rect 5442 6644 5448 6656
rect 5123 6616 5448 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 7098 6644 7104 6656
rect 6411 6616 7104 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 9232 6644 9260 6684
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 10873 6715 10931 6721
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 11146 6712 11152 6724
rect 10919 6684 11152 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 7515 6616 9260 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 12176 6644 12204 6752
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 15194 6780 15200 6792
rect 13127 6752 15200 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 12526 6712 12532 6724
rect 12308 6684 12532 6712
rect 12308 6672 12314 6684
rect 12526 6672 12532 6684
rect 12584 6672 12590 6724
rect 13906 6672 13912 6724
rect 13964 6712 13970 6724
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 13964 6684 14381 6712
rect 13964 6672 13970 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 14553 6715 14611 6721
rect 14553 6681 14565 6715
rect 14599 6712 14611 6715
rect 14918 6712 14924 6724
rect 14599 6684 14924 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 14918 6672 14924 6684
rect 14976 6672 14982 6724
rect 15654 6672 15660 6724
rect 15712 6712 15718 6724
rect 16114 6712 16120 6724
rect 15712 6684 16120 6712
rect 15712 6672 15718 6684
rect 16114 6672 16120 6684
rect 16172 6712 16178 6724
rect 16408 6712 16436 6743
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 16724 6752 17448 6780
rect 16724 6740 16730 6752
rect 16172 6684 16436 6712
rect 16172 6672 16178 6684
rect 16758 6672 16764 6724
rect 16816 6672 16822 6724
rect 17420 6712 17448 6752
rect 17494 6740 17500 6792
rect 17552 6740 17558 6792
rect 17604 6752 18644 6780
rect 17604 6712 17632 6752
rect 18230 6712 18236 6724
rect 17420 6684 17632 6712
rect 17926 6684 18236 6712
rect 9364 6616 12204 6644
rect 9364 6604 9370 6616
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13354 6644 13360 6656
rect 12676 6616 13360 6644
rect 12676 6604 12682 6616
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 14274 6644 14280 6656
rect 13771 6616 14280 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 15010 6604 15016 6656
rect 15068 6604 15074 6656
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 15381 6647 15439 6653
rect 15381 6644 15393 6647
rect 15344 6616 15393 6644
rect 15344 6604 15350 6616
rect 15381 6613 15393 6616
rect 15427 6613 15439 6647
rect 15381 6607 15439 6613
rect 15470 6604 15476 6656
rect 15528 6604 15534 6656
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 17926 6644 17954 6684
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 18616 6712 18644 6752
rect 19794 6740 19800 6792
rect 19852 6740 19858 6792
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 20916 6752 22661 6780
rect 18616 6684 19564 6712
rect 17644 6616 17954 6644
rect 17644 6604 17650 6616
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 18564 6616 19441 6644
rect 18564 6604 18570 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19536 6644 19564 6684
rect 20070 6672 20076 6724
rect 20128 6712 20134 6724
rect 20916 6712 20944 6752
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 24670 6740 24676 6792
rect 24728 6740 24734 6792
rect 20128 6684 20944 6712
rect 20128 6672 20134 6684
rect 21910 6672 21916 6724
rect 21968 6672 21974 6724
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 25038 6712 25044 6724
rect 23891 6684 25044 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 19536 6616 19901 6644
rect 19429 6607 19487 6613
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 934 6400 940 6452
rect 992 6440 998 6452
rect 3142 6440 3148 6452
rect 992 6412 3148 6440
rect 992 6400 998 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3375 6443 3433 6449
rect 3375 6409 3387 6443
rect 3421 6440 3433 6443
rect 3421 6412 7788 6440
rect 3421 6409 3433 6412
rect 3375 6403 3433 6409
rect 4709 6375 4767 6381
rect 4709 6341 4721 6375
rect 4755 6372 4767 6375
rect 5166 6372 5172 6384
rect 4755 6344 5172 6372
rect 4755 6341 4767 6344
rect 4709 6335 4767 6341
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 5258 6332 5264 6384
rect 5316 6372 5322 6384
rect 7650 6372 7656 6384
rect 5316 6344 7656 6372
rect 5316 6332 5322 6344
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 1627 6276 5365 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 5353 6273 5365 6276
rect 5399 6304 5411 6307
rect 5399 6276 7144 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 474 6196 480 6248
rect 532 6236 538 6248
rect 1857 6239 1915 6245
rect 1857 6236 1869 6239
rect 532 6208 1869 6236
rect 532 6196 538 6208
rect 1857 6205 1869 6208
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 2314 6236 2320 6248
rect 2179 6208 2320 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 1872 6100 1900 6199
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3878 6236 3884 6248
rect 3200 6208 3884 6236
rect 3200 6196 3206 6208
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4338 6196 4344 6248
rect 4396 6196 4402 6248
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 4982 6236 4988 6248
rect 4856 6208 4988 6236
rect 4856 6196 4862 6208
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 6730 6236 6736 6248
rect 6595 6208 6736 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 5997 6171 6055 6177
rect 2740 6140 4844 6168
rect 2740 6128 2746 6140
rect 4816 6112 4844 6140
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 7006 6168 7012 6180
rect 6043 6140 7012 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 7116 6168 7144 6276
rect 7190 6264 7196 6316
rect 7248 6264 7254 6316
rect 7760 6236 7788 6412
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 11149 6443 11207 6449
rect 11149 6440 11161 6443
rect 8812 6412 11161 6440
rect 8812 6400 8818 6412
rect 11149 6409 11161 6412
rect 11195 6440 11207 6443
rect 11330 6440 11336 6452
rect 11195 6412 11336 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 12805 6443 12863 6449
rect 12805 6440 12817 6443
rect 12084 6412 12817 6440
rect 7837 6375 7895 6381
rect 7837 6341 7849 6375
rect 7883 6372 7895 6375
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 7883 6344 9689 6372
rect 7883 6341 7895 6344
rect 7837 6335 7895 6341
rect 9677 6341 9689 6344
rect 9723 6341 9735 6375
rect 11606 6372 11612 6384
rect 10902 6344 11612 6372
rect 9677 6335 9735 6341
rect 11606 6332 11612 6344
rect 11664 6372 11670 6384
rect 11974 6372 11980 6384
rect 11664 6344 11980 6372
rect 11664 6332 11670 6344
rect 11974 6332 11980 6344
rect 12032 6372 12038 6384
rect 12084 6372 12112 6412
rect 12805 6409 12817 6412
rect 12851 6440 12863 6443
rect 13906 6440 13912 6452
rect 12851 6412 13912 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 14826 6440 14832 6452
rect 14056 6412 14832 6440
rect 14056 6400 14062 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15068 6412 16037 6440
rect 15068 6400 15074 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 17313 6443 17371 6449
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 17770 6440 17776 6452
rect 17359 6412 17776 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 20438 6440 20444 6452
rect 18248 6412 20444 6440
rect 12032 6344 12112 6372
rect 12032 6332 12038 6344
rect 12526 6332 12532 6384
rect 12584 6372 12590 6384
rect 13081 6375 13139 6381
rect 13081 6372 13093 6375
rect 12584 6344 13093 6372
rect 12584 6332 12590 6344
rect 13081 6341 13093 6344
rect 13127 6372 13139 6375
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13127 6344 13645 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 13633 6335 13691 6341
rect 14366 6332 14372 6384
rect 14424 6372 14430 6384
rect 15286 6372 15292 6384
rect 14424 6344 15292 6372
rect 14424 6332 14430 6344
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 15470 6332 15476 6384
rect 15528 6372 15534 6384
rect 15933 6375 15991 6381
rect 15933 6372 15945 6375
rect 15528 6344 15945 6372
rect 15528 6332 15534 6344
rect 15933 6341 15945 6344
rect 15979 6372 15991 6375
rect 16482 6372 16488 6384
rect 15979 6344 16488 6372
rect 15979 6341 15991 6344
rect 15933 6335 15991 6341
rect 16482 6332 16488 6344
rect 16540 6332 16546 6384
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 9214 6304 9220 6316
rect 8343 6276 9220 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 13538 6304 13544 6316
rect 12069 6267 12127 6273
rect 12912 6276 13544 6304
rect 9306 6236 9312 6248
rect 7760 6208 9312 6236
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9398 6196 9404 6248
rect 9456 6196 9462 6248
rect 11238 6236 11244 6248
rect 9508 6208 11244 6236
rect 9508 6168 9536 6208
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12084 6236 12112 6267
rect 11848 6208 12112 6236
rect 11848 6196 11854 6208
rect 12158 6196 12164 6248
rect 12216 6196 12222 6248
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 12912 6177 12940 6276
rect 13538 6264 13544 6276
rect 13596 6304 13602 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13596 6276 13737 6304
rect 13596 6264 13602 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14332 6276 14473 6304
rect 14332 6264 14338 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14608 6276 16252 6304
rect 14608 6264 14614 6276
rect 13814 6236 13820 6248
rect 13188 6208 13820 6236
rect 12897 6171 12955 6177
rect 12897 6168 12909 6171
rect 7116 6140 9536 6168
rect 11624 6140 12909 6168
rect 4154 6100 4160 6112
rect 1872 6072 4160 6100
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 4798 6060 4804 6112
rect 4856 6060 4862 6112
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 6730 6100 6736 6112
rect 6503 6072 6736 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 8570 6100 8576 6112
rect 6880 6072 8576 6100
rect 6880 6060 6886 6072
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 8938 6060 8944 6112
rect 8996 6060 9002 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 11624 6100 11652 6140
rect 12897 6137 12909 6140
rect 12943 6137 12955 6171
rect 12897 6131 12955 6137
rect 9180 6072 11652 6100
rect 11701 6103 11759 6109
rect 9180 6060 9186 6072
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 11974 6100 11980 6112
rect 11747 6072 11980 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 13188 6100 13216 6208
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 15194 6236 15200 6248
rect 13955 6208 15200 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 15838 6236 15844 6248
rect 15620 6208 15844 6236
rect 15620 6196 15626 6208
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 16114 6196 16120 6248
rect 16172 6196 16178 6248
rect 13265 6171 13323 6177
rect 13265 6137 13277 6171
rect 13311 6168 13323 6171
rect 15930 6168 15936 6180
rect 13311 6140 15936 6168
rect 13311 6137 13323 6140
rect 13265 6131 13323 6137
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 16224 6168 16252 6276
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 18248 6313 18276 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 21545 6443 21603 6449
rect 21545 6409 21557 6443
rect 21591 6440 21603 6443
rect 21726 6440 21732 6452
rect 21591 6412 21732 6440
rect 21591 6409 21603 6412
rect 21545 6403 21603 6409
rect 21726 6400 21732 6412
rect 21784 6400 21790 6452
rect 19242 6332 19248 6384
rect 19300 6332 19306 6384
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16448 6276 17233 6304
rect 16448 6264 16454 6276
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 20254 6264 20260 6316
rect 20312 6304 20318 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20312 6276 20821 6304
rect 20312 6264 20318 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 23937 6307 23995 6313
rect 23937 6273 23949 6307
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 16758 6196 16764 6248
rect 16816 6236 16822 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 16816 6208 17417 6236
rect 16816 6196 16822 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17586 6196 17592 6248
rect 17644 6236 17650 6248
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 17644 6208 18521 6236
rect 17644 6196 17650 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 18509 6199 18567 6205
rect 19536 6208 20913 6236
rect 16224 6140 17356 6168
rect 12400 6072 13216 6100
rect 12400 6060 12406 6072
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 13412 6072 15117 6100
rect 13412 6060 13418 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 15562 6060 15568 6112
rect 15620 6060 15626 6112
rect 16853 6103 16911 6109
rect 16853 6069 16865 6103
rect 16899 6100 16911 6103
rect 17218 6100 17224 6112
rect 16899 6072 17224 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 17328 6100 17356 6140
rect 17678 6128 17684 6180
rect 17736 6168 17742 6180
rect 17736 6140 18368 6168
rect 17736 6128 17742 6140
rect 17957 6103 18015 6109
rect 17957 6100 17969 6103
rect 17328 6072 17969 6100
rect 17957 6069 17969 6072
rect 18003 6100 18015 6103
rect 18230 6100 18236 6112
rect 18003 6072 18236 6100
rect 18003 6069 18015 6072
rect 17957 6063 18015 6069
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 18340 6100 18368 6140
rect 19536 6100 19564 6208
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 20901 6199 20959 6205
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6205 21051 6239
rect 20993 6199 21051 6205
rect 19702 6128 19708 6180
rect 19760 6168 19766 6180
rect 21008 6168 21036 6199
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 21784 6208 22477 6236
rect 21784 6196 21790 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 19760 6140 21036 6168
rect 19760 6128 19766 6140
rect 18340 6072 19564 6100
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 19981 6103 20039 6109
rect 19981 6100 19993 6103
rect 19668 6072 19993 6100
rect 19668 6060 19674 6072
rect 19981 6069 19993 6072
rect 20027 6069 20039 6103
rect 19981 6063 20039 6069
rect 20254 6060 20260 6112
rect 20312 6060 20318 6112
rect 20441 6103 20499 6109
rect 20441 6069 20453 6103
rect 20487 6100 20499 6103
rect 20530 6100 20536 6112
rect 20487 6072 20536 6100
rect 20487 6069 20499 6072
rect 20441 6063 20499 6069
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 20622 6060 20628 6112
rect 20680 6100 20686 6112
rect 23952 6100 23980 6267
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 20680 6072 23980 6100
rect 20680 6060 20686 6072
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 2682 5896 2688 5908
rect 1627 5868 2688 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 4617 5899 4675 5905
rect 4617 5896 4629 5899
rect 2832 5868 4629 5896
rect 2832 5856 2838 5868
rect 4617 5865 4629 5868
rect 4663 5865 4675 5899
rect 6822 5896 6828 5908
rect 4617 5859 4675 5865
rect 4724 5868 6828 5896
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4724 5828 4752 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 7248 5868 8585 5896
rect 7248 5856 7254 5868
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 8573 5859 8631 5865
rect 9122 5856 9128 5908
rect 9180 5856 9186 5908
rect 10045 5899 10103 5905
rect 10045 5865 10057 5899
rect 10091 5896 10103 5899
rect 11054 5896 11060 5908
rect 10091 5868 11060 5896
rect 10091 5865 10103 5868
rect 10045 5859 10103 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 11204 5868 12357 5896
rect 11204 5856 11210 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 12676 5868 12725 5896
rect 12676 5856 12682 5868
rect 12713 5865 12725 5868
rect 12759 5896 12771 5899
rect 13538 5896 13544 5908
rect 12759 5868 13544 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 13780 5868 17356 5896
rect 13780 5856 13786 5868
rect 4212 5800 4752 5828
rect 4212 5788 4218 5800
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 7282 5828 7288 5840
rect 4856 5800 7288 5828
rect 4856 5788 4862 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 7469 5831 7527 5837
rect 7469 5797 7481 5831
rect 7515 5828 7527 5831
rect 10505 5831 10563 5837
rect 7515 5800 10456 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 7650 5760 7656 5772
rect 2915 5732 7656 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 7800 5732 9904 5760
rect 7800 5720 7806 5732
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2406 5692 2412 5704
rect 1995 5664 2412 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2547 5664 2605 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2130 5584 2136 5636
rect 2188 5584 2194 5636
rect 2608 5624 2636 5655
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3844 5664 3985 5692
rect 3844 5652 3850 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 5031 5664 5089 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 5077 5661 5089 5664
rect 5123 5692 5135 5695
rect 5166 5692 5172 5704
rect 5123 5664 5172 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 4154 5624 4160 5636
rect 2608 5596 4160 5624
rect 4154 5584 4160 5596
rect 4212 5624 4218 5636
rect 4614 5624 4620 5636
rect 4212 5596 4620 5624
rect 4212 5584 4218 5596
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 6840 5624 6868 5655
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7616 5664 7941 5692
rect 7616 5652 7622 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 8996 5664 9413 5692
rect 8996 5652 9002 5664
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9582 5624 9588 5636
rect 6840 5596 9588 5624
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 3602 5516 3608 5568
rect 3660 5556 3666 5568
rect 3786 5556 3792 5568
rect 3660 5528 3792 5556
rect 3660 5516 3666 5528
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 6362 5516 6368 5568
rect 6420 5516 6426 5568
rect 9876 5556 9904 5732
rect 10428 5692 10456 5800
rect 10505 5797 10517 5831
rect 10551 5828 10563 5831
rect 12802 5828 12808 5840
rect 10551 5800 12808 5828
rect 10551 5797 10563 5800
rect 10505 5791 10563 5797
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 14277 5831 14335 5837
rect 14277 5797 14289 5831
rect 14323 5828 14335 5831
rect 14366 5828 14372 5840
rect 14323 5800 14372 5828
rect 14323 5797 14335 5800
rect 14277 5791 14335 5797
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 15194 5828 15200 5840
rect 14792 5800 15200 5828
rect 14792 5788 14798 5800
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 17328 5828 17356 5868
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 18877 5899 18935 5905
rect 18877 5896 18889 5899
rect 17460 5868 18889 5896
rect 17460 5856 17466 5868
rect 18877 5865 18889 5868
rect 18923 5865 18935 5899
rect 18877 5859 18935 5865
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 20254 5896 20260 5908
rect 19300 5868 20260 5896
rect 19300 5856 19306 5868
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 23290 5896 23296 5908
rect 21692 5868 23296 5896
rect 21692 5856 21698 5868
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 17328 5800 18276 5828
rect 10594 5720 10600 5772
rect 10652 5760 10658 5772
rect 11057 5763 11115 5769
rect 11057 5760 11069 5763
rect 10652 5732 11069 5760
rect 10652 5720 10658 5732
rect 11057 5729 11069 5732
rect 11103 5729 11115 5763
rect 17586 5760 17592 5772
rect 11057 5723 11115 5729
rect 11164 5732 11836 5760
rect 11164 5692 11192 5732
rect 10428 5664 11192 5692
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11808 5692 11836 5732
rect 13004 5732 17592 5760
rect 13004 5692 13032 5732
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 11808 5664 13032 5692
rect 13081 5695 13139 5701
rect 11701 5655 11759 5661
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13354 5692 13360 5704
rect 13127 5664 13360 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 11716 5624 11744 5655
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 14734 5652 14740 5704
rect 14792 5652 14798 5704
rect 16022 5652 16028 5704
rect 16080 5652 16086 5704
rect 18138 5692 18144 5704
rect 17434 5664 18144 5692
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18248 5701 18276 5800
rect 18690 5788 18696 5840
rect 18748 5828 18754 5840
rect 18748 5800 21864 5828
rect 18748 5788 18754 5800
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19889 5763 19947 5769
rect 19889 5760 19901 5763
rect 19392 5732 19901 5760
rect 19392 5720 19398 5732
rect 19889 5729 19901 5732
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 21729 5763 21787 5769
rect 21729 5760 21741 5763
rect 20588 5732 21741 5760
rect 20588 5720 20594 5732
rect 21729 5729 21741 5732
rect 21775 5729 21787 5763
rect 21729 5723 21787 5729
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 20864 5664 21281 5692
rect 20864 5652 20870 5664
rect 21269 5661 21281 5664
rect 21315 5661 21327 5695
rect 21836 5692 21864 5800
rect 23477 5763 23535 5769
rect 23477 5729 23489 5763
rect 23523 5760 23535 5763
rect 23566 5760 23572 5772
rect 23523 5732 23572 5760
rect 23523 5729 23535 5732
rect 23477 5723 23535 5729
rect 23566 5720 23572 5732
rect 23624 5720 23630 5772
rect 24026 5720 24032 5772
rect 24084 5760 24090 5772
rect 25041 5763 25099 5769
rect 25041 5760 25053 5763
rect 24084 5732 25053 5760
rect 24084 5720 24090 5732
rect 25041 5729 25053 5732
rect 25087 5729 25099 5763
rect 25041 5723 25099 5729
rect 25225 5763 25283 5769
rect 25225 5729 25237 5763
rect 25271 5760 25283 5763
rect 25314 5760 25320 5772
rect 25271 5732 25320 5760
rect 25271 5729 25283 5732
rect 25225 5723 25283 5729
rect 25314 5720 25320 5732
rect 25372 5720 25378 5772
rect 22830 5692 22836 5704
rect 21836 5664 22836 5692
rect 21269 5655 21327 5661
rect 22830 5652 22836 5664
rect 22888 5652 22894 5704
rect 23201 5695 23259 5701
rect 23201 5661 23213 5695
rect 23247 5692 23259 5695
rect 24486 5692 24492 5704
rect 23247 5664 24492 5692
rect 23247 5661 23259 5664
rect 23201 5655 23259 5661
rect 24486 5652 24492 5664
rect 24544 5652 24550 5704
rect 10836 5596 11744 5624
rect 10836 5584 10842 5596
rect 15102 5584 15108 5636
rect 15160 5624 15166 5636
rect 16301 5627 16359 5633
rect 16301 5624 16313 5627
rect 15160 5596 16313 5624
rect 15160 5584 15166 5596
rect 16301 5593 16313 5596
rect 16347 5593 16359 5627
rect 19978 5624 19984 5636
rect 16301 5587 16359 5593
rect 17696 5596 19984 5624
rect 10873 5559 10931 5565
rect 10873 5556 10885 5559
rect 9876 5528 10885 5556
rect 10873 5525 10885 5528
rect 10919 5525 10931 5559
rect 10873 5519 10931 5525
rect 10962 5516 10968 5568
rect 11020 5516 11026 5568
rect 13354 5516 13360 5568
rect 13412 5556 13418 5568
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 13412 5528 13737 5556
rect 13412 5516 13418 5528
rect 13725 5525 13737 5528
rect 13771 5525 13783 5559
rect 13725 5519 13783 5525
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14458 5556 14464 5568
rect 13964 5528 14464 5556
rect 13964 5516 13970 5528
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 14967 5559 15025 5565
rect 14967 5525 14979 5559
rect 15013 5556 15025 5559
rect 17696 5556 17724 5596
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 20714 5584 20720 5636
rect 20772 5624 20778 5636
rect 24397 5627 24455 5633
rect 24397 5624 24409 5627
rect 20772 5596 24409 5624
rect 20772 5584 20778 5596
rect 24397 5593 24409 5596
rect 24443 5624 24455 5627
rect 24949 5627 25007 5633
rect 24949 5624 24961 5627
rect 24443 5596 24961 5624
rect 24443 5593 24455 5596
rect 24397 5587 24455 5593
rect 24949 5593 24961 5596
rect 24995 5593 25007 5627
rect 24949 5587 25007 5593
rect 15013 5528 17724 5556
rect 15013 5525 15025 5528
rect 14967 5519 15025 5525
rect 17770 5516 17776 5568
rect 17828 5516 17834 5568
rect 20438 5516 20444 5568
rect 20496 5556 20502 5568
rect 22002 5556 22008 5568
rect 20496 5528 22008 5556
rect 20496 5516 20502 5528
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 24578 5516 24584 5568
rect 24636 5516 24642 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 3970 5352 3976 5364
rect 2271 5324 3976 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 5074 5312 5080 5364
rect 5132 5312 5138 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 7374 5352 7380 5364
rect 5408 5324 7380 5352
rect 5408 5312 5414 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7708 5324 7849 5352
rect 7708 5312 7714 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 15102 5352 15108 5364
rect 11195 5324 15108 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 15930 5312 15936 5364
rect 15988 5312 15994 5364
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 16540 5324 16865 5352
rect 16540 5312 16546 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 16853 5315 16911 5321
rect 17126 5312 17132 5364
rect 17184 5312 17190 5364
rect 19610 5312 19616 5364
rect 19668 5352 19674 5364
rect 21177 5355 21235 5361
rect 21177 5352 21189 5355
rect 19668 5324 21189 5352
rect 19668 5312 19674 5324
rect 21177 5321 21189 5324
rect 21223 5321 21235 5355
rect 21177 5315 21235 5321
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22738 5352 22744 5364
rect 22152 5324 22744 5352
rect 22152 5312 22158 5324
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 12158 5284 12164 5296
rect 4172 5256 12164 5284
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 3602 5216 3608 5228
rect 2731 5188 3608 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 1596 5148 1624 5179
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4172 5225 4200 5256
rect 12158 5244 12164 5256
rect 12216 5244 12222 5296
rect 13354 5244 13360 5296
rect 13412 5244 13418 5296
rect 16942 5284 16948 5296
rect 14752 5256 16948 5284
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 6086 5216 6092 5228
rect 5399 5188 6092 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 7156 5188 7205 5216
rect 7156 5176 7162 5188
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 9306 5216 9312 5228
rect 8343 5188 9312 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9950 5216 9956 5228
rect 9447 5188 9956 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10091 5188 10517 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 11606 5176 11612 5228
rect 11664 5176 11670 5228
rect 11974 5176 11980 5228
rect 12032 5176 12038 5228
rect 14458 5176 14464 5228
rect 14516 5176 14522 5228
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 1596 5120 3341 5148
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 3896 5080 3924 5111
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 6549 5151 6607 5157
rect 4764 5120 6500 5148
rect 4764 5108 4770 5120
rect 6086 5080 6092 5092
rect 3896 5052 6092 5080
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 6472 5080 6500 5120
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 12250 5148 12256 5160
rect 6595 5120 12256 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 12986 5148 12992 5160
rect 12768 5120 12992 5148
rect 12768 5108 12774 5120
rect 12986 5108 12992 5120
rect 13044 5148 13050 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 13044 5120 13093 5148
rect 13044 5108 13050 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 14642 5148 14648 5160
rect 13081 5111 13139 5117
rect 13188 5120 14648 5148
rect 13188 5080 13216 5120
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 6472 5052 13216 5080
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 14752 5080 14780 5256
rect 16942 5244 16948 5256
rect 17000 5284 17006 5296
rect 17770 5284 17776 5296
rect 17000 5256 17776 5284
rect 17000 5244 17006 5256
rect 17770 5244 17776 5256
rect 17828 5244 17834 5296
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15344 5188 15853 5216
rect 15344 5176 15350 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 16356 5188 17417 5216
rect 16356 5176 16362 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 14424 5052 14780 5080
rect 14844 5120 16037 5148
rect 14424 5040 14430 5052
rect 14844 5024 14872 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 18322 5108 18328 5160
rect 18380 5108 18386 5160
rect 14918 5040 14924 5092
rect 14976 5080 14982 5092
rect 19260 5080 19288 5179
rect 21174 5176 21180 5228
rect 21232 5216 21238 5228
rect 21361 5219 21419 5225
rect 21361 5216 21373 5219
rect 21232 5188 21373 5216
rect 21232 5176 21238 5188
rect 21361 5185 21373 5188
rect 21407 5185 21419 5219
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21361 5179 21419 5185
rect 21468 5188 22017 5216
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5117 19763 5151
rect 19705 5111 19763 5117
rect 14976 5052 19288 5080
rect 14976 5040 14982 5052
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4338 5012 4344 5024
rect 4212 4984 4344 5012
rect 4212 4972 4218 4984
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 5997 5015 6055 5021
rect 5997 4981 6009 5015
rect 6043 5012 6055 5015
rect 8846 5012 8852 5024
rect 6043 4984 8852 5012
rect 6043 4981 6055 4984
rect 5997 4975 6055 4981
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 8938 4972 8944 5024
rect 8996 4972 9002 5024
rect 10318 4972 10324 5024
rect 10376 5012 10382 5024
rect 11606 5012 11612 5024
rect 10376 4984 11612 5012
rect 10376 4972 10382 4984
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12621 5015 12679 5021
rect 12621 4981 12633 5015
rect 12667 5012 12679 5015
rect 12802 5012 12808 5024
rect 12667 4984 12808 5012
rect 12667 4981 12679 4984
rect 12621 4975 12679 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 13446 5012 13452 5024
rect 13044 4984 13452 5012
rect 13044 4972 13050 4984
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 14826 4972 14832 5024
rect 14884 4972 14890 5024
rect 15286 4972 15292 5024
rect 15344 4972 15350 5024
rect 15470 4972 15476 5024
rect 15528 4972 15534 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17862 5012 17868 5024
rect 17460 4984 17868 5012
rect 17460 4972 17466 4984
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 19720 5012 19748 5111
rect 19794 5108 19800 5160
rect 19852 5148 19858 5160
rect 21468 5148 21496 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 23934 5176 23940 5228
rect 23992 5176 23998 5228
rect 19852 5120 21496 5148
rect 19852 5108 19858 5120
rect 21542 5108 21548 5160
rect 21600 5148 21606 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 21600 5120 22477 5148
rect 21600 5108 21606 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 18656 4984 19748 5012
rect 18656 4972 18662 4984
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 1872 4780 7604 4808
rect 1872 4681 1900 4780
rect 7576 4740 7604 4780
rect 7650 4768 7656 4820
rect 7708 4768 7714 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 8536 4780 8585 4808
rect 8536 4768 8542 4780
rect 8573 4777 8585 4780
rect 8619 4777 8631 4811
rect 8573 4771 8631 4777
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 9088 4780 9137 4808
rect 9088 4768 9094 4780
rect 9125 4777 9137 4780
rect 9171 4777 9183 4811
rect 9125 4771 9183 4777
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 15470 4808 15476 4820
rect 9364 4780 15476 4808
rect 9364 4768 9370 4780
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 15988 4780 16528 4808
rect 15988 4768 15994 4780
rect 16500 4752 16528 4780
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 19886 4808 19892 4820
rect 17828 4780 19892 4808
rect 17828 4768 17834 4780
rect 19886 4768 19892 4780
rect 19944 4808 19950 4820
rect 22189 4811 22247 4817
rect 22189 4808 22201 4811
rect 19944 4780 22201 4808
rect 19944 4768 19950 4780
rect 22189 4777 22201 4780
rect 22235 4777 22247 4811
rect 22189 4771 22247 4777
rect 14550 4740 14556 4752
rect 7576 4712 9674 4740
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 9398 4672 9404 4684
rect 5123 4644 9404 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9646 4672 9674 4712
rect 9784 4712 14556 4740
rect 9784 4672 9812 4712
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 14645 4743 14703 4749
rect 14645 4709 14657 4743
rect 14691 4740 14703 4743
rect 14918 4740 14924 4752
rect 14691 4712 14924 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 16482 4700 16488 4752
rect 16540 4740 16546 4752
rect 19061 4743 19119 4749
rect 19061 4740 19073 4743
rect 16540 4712 19073 4740
rect 16540 4700 16546 4712
rect 19061 4709 19073 4712
rect 19107 4740 19119 4743
rect 19702 4740 19708 4752
rect 19107 4712 19708 4740
rect 19107 4709 19119 4712
rect 19061 4703 19119 4709
rect 19702 4700 19708 4712
rect 19760 4740 19766 4752
rect 19760 4712 20576 4740
rect 19760 4700 19766 4712
rect 14826 4672 14832 4684
rect 9646 4644 9812 4672
rect 12406 4644 14832 4672
rect 1026 4564 1032 4616
rect 1084 4604 1090 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1084 4576 1593 4604
rect 1084 4564 1090 4576
rect 1581 4573 1593 4576
rect 1627 4604 1639 4607
rect 1762 4604 1768 4616
rect 1627 4576 1768 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 2924 4576 3249 4604
rect 2924 4564 2930 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3476 4576 3985 4604
rect 3476 4564 3482 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7147 4576 7941 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 7929 4573 7941 4576
rect 7975 4604 7987 4607
rect 8386 4604 8392 4616
rect 7975 4576 8392 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 9030 4604 9036 4616
rect 8536 4576 9036 4604
rect 8536 4564 8542 4576
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 9306 4564 9312 4616
rect 9364 4564 9370 4616
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 12406 4604 12434 4644
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 16022 4672 16028 4684
rect 15151 4644 16028 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 16172 4644 16865 4672
rect 16172 4632 16178 4644
rect 16853 4641 16865 4644
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 17862 4632 17868 4684
rect 17920 4672 17926 4684
rect 20257 4675 20315 4681
rect 20257 4672 20269 4675
rect 17920 4644 20269 4672
rect 17920 4632 17926 4644
rect 20257 4641 20269 4644
rect 20303 4641 20315 4675
rect 20257 4635 20315 4641
rect 12023 4576 12434 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 3344 4508 5304 4536
rect 2866 4428 2872 4480
rect 2924 4428 2930 4480
rect 3344 4477 3372 4508
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4437 3387 4471
rect 3329 4431 3387 4437
rect 4062 4428 4068 4480
rect 4120 4468 4126 4480
rect 4430 4468 4436 4480
rect 4120 4440 4436 4468
rect 4120 4428 4126 4440
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 4617 4471 4675 4477
rect 4617 4437 4629 4471
rect 4663 4468 4675 4471
rect 4798 4468 4804 4480
rect 4663 4440 4804 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5276 4468 5304 4508
rect 5350 4496 5356 4548
rect 5408 4496 5414 4548
rect 6578 4508 8294 4536
rect 6638 4468 6644 4480
rect 5276 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7469 4471 7527 4477
rect 7469 4437 7481 4471
rect 7515 4468 7527 4471
rect 7650 4468 7656 4480
rect 7515 4440 7656 4468
rect 7515 4437 7527 4440
rect 7469 4431 7527 4437
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 8266 4468 8294 4508
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 10413 4539 10471 4545
rect 10413 4536 10425 4539
rect 9272 4508 10425 4536
rect 9272 4496 9278 4508
rect 10413 4505 10425 4508
rect 10459 4505 10471 4539
rect 10888 4536 10916 4567
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 12860 4576 13093 4604
rect 12860 4564 12866 4576
rect 13081 4573 13093 4576
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13771 4576 14596 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 12621 4539 12679 4545
rect 12621 4536 12633 4539
rect 10888 4508 12633 4536
rect 10413 4499 10471 4505
rect 12621 4505 12633 4508
rect 12667 4505 12679 4539
rect 12621 4499 12679 4505
rect 14461 4539 14519 4545
rect 14461 4505 14473 4539
rect 14507 4505 14519 4539
rect 14568 4536 14596 4576
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 16684 4576 17325 4604
rect 15381 4539 15439 4545
rect 15381 4536 15393 4539
rect 14568 4508 15393 4536
rect 14461 4499 14519 4505
rect 15381 4505 15393 4508
rect 15427 4505 15439 4539
rect 15381 4499 15439 4505
rect 10318 4468 10324 4480
rect 8266 4440 10324 4468
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 10560 4440 11529 4468
rect 10560 4428 10566 4440
rect 11517 4437 11529 4440
rect 11563 4437 11575 4471
rect 11517 4431 11575 4437
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14476 4468 14504 4499
rect 14642 4468 14648 4480
rect 13780 4440 14648 4468
rect 13780 4428 13786 4440
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 14734 4428 14740 4480
rect 14792 4468 14798 4480
rect 16684 4468 16712 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 20070 4604 20076 4616
rect 19484 4576 20076 4604
rect 19484 4564 19490 4576
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 18414 4496 18420 4548
rect 18472 4496 18478 4548
rect 19242 4496 19248 4548
rect 19300 4536 19306 4548
rect 19705 4539 19763 4545
rect 19705 4536 19717 4539
rect 19300 4508 19717 4536
rect 19300 4496 19306 4508
rect 19705 4505 19717 4508
rect 19751 4505 19763 4539
rect 20272 4536 20300 4635
rect 20438 4632 20444 4684
rect 20496 4632 20502 4684
rect 20548 4672 20576 4712
rect 20806 4672 20812 4684
rect 20548 4644 20812 4672
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 21082 4632 21088 4684
rect 21140 4672 21146 4684
rect 23109 4675 23167 4681
rect 23109 4672 23121 4675
rect 21140 4644 23121 4672
rect 21140 4632 21146 4644
rect 23109 4641 23121 4644
rect 23155 4641 23167 4675
rect 23109 4635 23167 4641
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 24578 4564 24584 4616
rect 24636 4564 24642 4616
rect 20717 4539 20775 4545
rect 20717 4536 20729 4539
rect 20272 4508 20729 4536
rect 19705 4499 19763 4505
rect 20717 4505 20729 4508
rect 20763 4505 20775 4539
rect 20717 4499 20775 4505
rect 20806 4496 20812 4548
rect 20864 4536 20870 4548
rect 21174 4536 21180 4548
rect 20864 4508 21180 4536
rect 20864 4496 20870 4508
rect 21174 4496 21180 4508
rect 21232 4496 21238 4548
rect 22066 4508 22324 4536
rect 14792 4440 16712 4468
rect 14792 4428 14798 4440
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 22066 4468 22094 4508
rect 17368 4440 22094 4468
rect 22296 4468 22324 4508
rect 25225 4471 25283 4477
rect 25225 4468 25237 4471
rect 22296 4440 25237 4468
rect 17368 4428 17374 4440
rect 25225 4437 25237 4440
rect 25271 4437 25283 4471
rect 25225 4431 25283 4437
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 3234 4264 3240 4276
rect 2915 4236 3240 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 5408 4236 5457 4264
rect 5408 4224 5414 4236
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5445 4227 5503 4233
rect 6086 4224 6092 4276
rect 6144 4264 6150 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6144 4236 6561 4264
rect 6144 4224 6150 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7650 4264 7656 4276
rect 7156 4236 7656 4264
rect 7156 4224 7162 4236
rect 7650 4224 7656 4236
rect 7708 4264 7714 4276
rect 7708 4236 9536 4264
rect 7708 4224 7714 4236
rect 2958 4196 2964 4208
rect 1596 4168 2964 4196
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1596 4137 1624 4168
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 8754 4196 8760 4208
rect 6748 4168 8760 4196
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1544 4100 1593 4128
rect 1544 4088 1550 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2823 4100 3065 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 3053 4097 3065 4100
rect 3099 4128 3111 4131
rect 3326 4128 3332 4140
rect 3099 4100 3332 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5626 4128 5632 4140
rect 5040 4100 5632 4128
rect 5040 4088 5046 4100
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 5902 4128 5908 4140
rect 5859 4100 5908 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 6748 4137 6776 4168
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 7064 4100 7205 4128
rect 7064 4088 7070 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 2406 4060 2412 4072
rect 1903 4032 2412 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 3510 4020 3516 4072
rect 3568 4020 3574 4072
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4060 3847 4063
rect 5258 4060 5264 4072
rect 3835 4032 5264 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 8312 4060 8340 4091
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 8996 4100 9413 4128
rect 8996 4088 9002 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9508 4128 9536 4236
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 14366 4264 14372 4276
rect 9824 4236 14372 4264
rect 9824 4224 9830 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 14458 4224 14464 4276
rect 14516 4264 14522 4276
rect 15838 4264 15844 4276
rect 14516 4236 15844 4264
rect 14516 4224 14522 4236
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 14274 4196 14280 4208
rect 9732 4168 14280 4196
rect 9732 4156 9738 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 15580 4196 15608 4236
rect 15838 4224 15844 4236
rect 15896 4264 15902 4276
rect 16022 4264 16028 4276
rect 15896 4236 16028 4264
rect 15896 4224 15902 4236
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 17126 4224 17132 4276
rect 17184 4264 17190 4276
rect 17405 4267 17463 4273
rect 17405 4264 17417 4267
rect 17184 4236 17417 4264
rect 17184 4224 17190 4236
rect 17405 4233 17417 4236
rect 17451 4233 17463 4267
rect 18782 4264 18788 4276
rect 17405 4227 17463 4233
rect 17972 4236 18788 4264
rect 15502 4168 15608 4196
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 17972 4196 18000 4236
rect 18782 4224 18788 4236
rect 18840 4264 18846 4276
rect 19242 4264 19248 4276
rect 18840 4236 19248 4264
rect 18840 4224 18846 4236
rect 19242 4224 19248 4236
rect 19300 4264 19306 4276
rect 24302 4264 24308 4276
rect 19300 4236 24308 4264
rect 19300 4224 19306 4236
rect 24302 4224 24308 4236
rect 24360 4224 24366 4276
rect 18506 4196 18512 4208
rect 15712 4168 16574 4196
rect 15712 4156 15718 4168
rect 10134 4128 10140 4140
rect 9508 4100 10140 4128
rect 9401 4091 9459 4097
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11020 4100 11529 4128
rect 11020 4088 11026 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 12158 4088 12164 4140
rect 12216 4088 12222 4140
rect 13354 4088 13360 4140
rect 13412 4088 13418 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13504 4100 14013 4128
rect 13504 4088 13510 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 16209 4131 16267 4137
rect 16209 4128 16221 4131
rect 14001 4091 14059 4097
rect 15488 4100 16221 4128
rect 10042 4060 10048 4072
rect 8312 4032 10048 4060
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 11882 4060 11888 4072
rect 10152 4032 11888 4060
rect 2958 3952 2964 4004
rect 3016 3992 3022 4004
rect 10152 3992 10180 4032
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13372 4032 14289 4060
rect 3016 3964 10180 3992
rect 11149 3995 11207 4001
rect 3016 3952 3022 3964
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 13372 3992 13400 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 15488 4060 15516 4100
rect 16209 4097 16221 4100
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 16390 4088 16396 4140
rect 16448 4088 16454 4140
rect 16546 4128 16574 4168
rect 17420 4168 18000 4196
rect 18248 4168 18512 4196
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 16546 4100 16773 4128
rect 16761 4097 16773 4100
rect 16807 4128 16819 4131
rect 17420 4128 17448 4168
rect 16807 4100 17448 4128
rect 17497 4131 17555 4137
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 18248 4128 18276 4168
rect 18506 4156 18512 4168
rect 18564 4156 18570 4208
rect 19886 4156 19892 4208
rect 19944 4196 19950 4208
rect 21358 4196 21364 4208
rect 19944 4168 21364 4196
rect 19944 4156 19950 4168
rect 21358 4156 21364 4168
rect 21416 4156 21422 4208
rect 17543 4100 18276 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 19610 4088 19616 4140
rect 19668 4088 19674 4140
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 21542 4128 21548 4140
rect 20312 4100 21548 4128
rect 20312 4088 20318 4100
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 22186 4088 22192 4140
rect 22244 4088 22250 4140
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 23566 4128 23572 4140
rect 22888 4100 23572 4128
rect 22888 4088 22894 4100
rect 23566 4088 23572 4100
rect 23624 4088 23630 4140
rect 23842 4088 23848 4140
rect 23900 4088 23906 4140
rect 23934 4088 23940 4140
rect 23992 4128 23998 4140
rect 24946 4128 24952 4140
rect 23992 4100 24952 4128
rect 23992 4088 23998 4100
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 17586 4060 17592 4072
rect 14700 4032 15516 4060
rect 15672 4032 17592 4060
rect 14700 4020 14706 4032
rect 11195 3964 13400 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4430 3924 4436 3936
rect 3844 3896 4436 3924
rect 3844 3884 3850 3896
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 5902 3884 5908 3936
rect 5960 3884 5966 3936
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6454 3924 6460 3936
rect 6227 3896 6460 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7800 3896 7849 3924
rect 7800 3884 7806 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 7837 3887 7895 3893
rect 8938 3884 8944 3936
rect 8996 3884 9002 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10045 3927 10103 3933
rect 10045 3924 10057 3927
rect 9732 3896 10057 3924
rect 9732 3884 9738 3896
rect 10045 3893 10057 3896
rect 10091 3893 10103 3927
rect 10045 3887 10103 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 10192 3896 11897 3924
rect 10192 3884 10198 3896
rect 11885 3893 11897 3896
rect 11931 3924 11943 3927
rect 12618 3924 12624 3936
rect 11931 3896 12624 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 15672 3924 15700 4032
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 18233 4063 18291 4069
rect 18233 4029 18245 4063
rect 18279 4029 18291 4063
rect 18233 4023 18291 4029
rect 12768 3896 15700 3924
rect 12768 3884 12774 3896
rect 15746 3884 15752 3936
rect 15804 3884 15810 3936
rect 16022 3884 16028 3936
rect 16080 3884 16086 3936
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 17037 3927 17095 3933
rect 17037 3924 17049 3927
rect 16816 3896 17049 3924
rect 16816 3884 16822 3896
rect 17037 3893 17049 3896
rect 17083 3893 17095 3927
rect 18248 3924 18276 4023
rect 18506 4020 18512 4072
rect 18564 4020 18570 4072
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 20346 4060 20352 4072
rect 19760 4032 20352 4060
rect 19760 4020 19766 4032
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 20625 4063 20683 4069
rect 20625 4029 20637 4063
rect 20671 4060 20683 4063
rect 20714 4060 20720 4072
rect 20671 4032 20720 4060
rect 20671 4029 20683 4032
rect 20625 4023 20683 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 20901 4063 20959 4069
rect 20901 4060 20913 4063
rect 20864 4032 20913 4060
rect 20864 4020 20870 4032
rect 20901 4029 20913 4032
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 21450 4020 21456 4072
rect 21508 4060 21514 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 21508 4032 22477 4060
rect 21508 4020 21514 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 21358 3952 21364 4004
rect 21416 3992 21422 4004
rect 24320 3992 24348 4023
rect 21416 3964 24348 3992
rect 21416 3952 21422 3964
rect 19702 3924 19708 3936
rect 18248 3896 19708 3924
rect 17037 3887 17095 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 19978 3884 19984 3936
rect 20036 3884 20042 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20346 3924 20352 3936
rect 20220 3896 20352 3924
rect 20220 3884 20226 3896
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 21634 3884 21640 3936
rect 21692 3924 21698 3936
rect 24946 3924 24952 3936
rect 21692 3896 24952 3924
rect 21692 3884 21698 3896
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2041 3723 2099 3729
rect 2041 3689 2053 3723
rect 2087 3720 2099 3723
rect 2087 3692 2774 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 2746 3652 2774 3692
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3786 3720 3792 3732
rect 3476 3692 3792 3720
rect 3476 3680 3482 3692
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 7006 3720 7012 3732
rect 4580 3692 7012 3720
rect 4580 3680 4586 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 7432 3692 9137 3720
rect 7432 3680 7438 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 10686 3720 10692 3732
rect 9125 3683 9183 3689
rect 9232 3692 10692 3720
rect 5718 3652 5724 3664
rect 2556 3624 2636 3652
rect 2746 3624 5724 3652
rect 2556 3612 2562 3624
rect 2608 3593 2636 3624
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 5994 3612 6000 3664
rect 6052 3652 6058 3664
rect 6365 3655 6423 3661
rect 6365 3652 6377 3655
rect 6052 3624 6377 3652
rect 6052 3612 6058 3624
rect 6365 3621 6377 3624
rect 6411 3652 6423 3655
rect 7098 3652 7104 3664
rect 6411 3624 7104 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 7098 3612 7104 3624
rect 7156 3612 7162 3664
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3553 2651 3587
rect 3234 3584 3240 3596
rect 2593 3547 2651 3553
rect 2746 3556 3240 3584
rect 658 3476 664 3528
rect 716 3516 722 3528
rect 1394 3516 1400 3528
rect 716 3488 1400 3516
rect 716 3476 722 3488
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1912 3488 1961 3516
rect 1912 3476 1918 3488
rect 1949 3485 1961 3488
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2746 3516 2774 3556
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 3786 3544 3792 3596
rect 3844 3584 3850 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 3844 3556 3985 3584
rect 3844 3544 3850 3556
rect 3973 3553 3985 3556
rect 4019 3584 4031 3587
rect 4338 3584 4344 3596
rect 4019 3556 4344 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 9232 3584 9260 3692
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 11974 3720 11980 3732
rect 11563 3692 11980 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 15930 3720 15936 3732
rect 12676 3692 15936 3720
rect 12676 3680 12682 3692
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 18322 3720 18328 3732
rect 17368 3692 18328 3720
rect 17368 3680 17374 3692
rect 18322 3680 18328 3692
rect 18380 3680 18386 3732
rect 23842 3720 23848 3732
rect 18800 3692 23848 3720
rect 16758 3652 16764 3664
rect 5184 3556 9260 3584
rect 9324 3624 16764 3652
rect 2096 3488 2774 3516
rect 2096 3476 2102 3488
rect 2866 3476 2872 3528
rect 2924 3476 2930 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 4154 3516 4160 3528
rect 3476 3488 4160 3516
rect 3476 3476 3482 3488
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 5184 3516 5212 3556
rect 4295 3488 5212 3516
rect 5261 3519 5319 3525
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 2958 3448 2964 3460
rect 1627 3420 2964 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 5276 3448 5304 3479
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 9324 3525 9352 3624
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 16942 3612 16948 3664
rect 17000 3652 17006 3664
rect 18414 3652 18420 3664
rect 17000 3624 18420 3652
rect 17000 3612 17006 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 12710 3584 12716 3596
rect 9784 3556 12716 3584
rect 9784 3525 9812 3556
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 18046 3544 18052 3596
rect 18104 3544 18110 3596
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3516 10931 3519
rect 12529 3519 12587 3525
rect 10919 3488 12434 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 3712 3420 5304 3448
rect 6549 3451 6607 3457
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 3712 3380 3740 3420
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 11698 3448 11704 3460
rect 6595 3420 11704 3448
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3448 11943 3451
rect 12066 3448 12072 3460
rect 11931 3420 12072 3448
rect 11931 3417 11943 3420
rect 11885 3411 11943 3417
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12406 3448 12434 3488
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 13446 3516 13452 3528
rect 12575 3488 13452 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 15746 3516 15752 3528
rect 15028 3488 15752 3516
rect 15028 3448 15056 3488
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 16206 3476 16212 3528
rect 16264 3476 16270 3528
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18690 3516 18696 3528
rect 18371 3488 18696 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 12406 3420 15056 3448
rect 15102 3408 15108 3460
rect 15160 3448 15166 3460
rect 18800 3448 18828 3692
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24210 3680 24216 3732
rect 24268 3680 24274 3732
rect 23290 3612 23296 3664
rect 23348 3612 23354 3664
rect 23658 3612 23664 3664
rect 23716 3612 23722 3664
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3584 19487 3587
rect 19702 3584 19708 3596
rect 19475 3556 19708 3584
rect 19475 3553 19487 3556
rect 19429 3547 19487 3553
rect 19702 3544 19708 3556
rect 19760 3584 19766 3596
rect 20438 3584 20444 3596
rect 19760 3556 20444 3584
rect 19760 3544 19766 3556
rect 20438 3544 20444 3556
rect 20496 3544 20502 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 22097 3587 22155 3593
rect 22097 3584 22109 3587
rect 20772 3556 22109 3584
rect 20772 3544 20778 3556
rect 22097 3553 22109 3556
rect 22143 3553 22155 3587
rect 22097 3547 22155 3553
rect 22554 3544 22560 3596
rect 22612 3584 22618 3596
rect 23477 3587 23535 3593
rect 23477 3584 23489 3587
rect 22612 3556 23489 3584
rect 22612 3544 22618 3556
rect 23308 3528 23336 3556
rect 23477 3553 23489 3556
rect 23523 3553 23535 3587
rect 23477 3547 23535 3553
rect 21174 3516 21180 3528
rect 20838 3488 21180 3516
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 21634 3476 21640 3528
rect 21692 3476 21698 3528
rect 23290 3476 23296 3528
rect 23348 3476 23354 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24486 3516 24492 3528
rect 24360 3488 24492 3516
rect 24360 3476 24366 3488
rect 24486 3476 24492 3488
rect 24544 3516 24550 3528
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24544 3488 24685 3516
rect 24544 3476 24550 3488
rect 24673 3485 24685 3488
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 15160 3420 18828 3448
rect 15160 3408 15166 3420
rect 19702 3408 19708 3460
rect 19760 3408 19766 3460
rect 21192 3448 21220 3476
rect 22002 3448 22008 3460
rect 21192 3420 22008 3448
rect 22002 3408 22008 3420
rect 22060 3448 22066 3460
rect 24210 3448 24216 3460
rect 22060 3420 24216 3448
rect 22060 3408 22066 3420
rect 24210 3408 24216 3420
rect 24268 3448 24274 3460
rect 25041 3451 25099 3457
rect 25041 3448 25053 3451
rect 24268 3420 25053 3448
rect 24268 3408 24274 3420
rect 25041 3417 25053 3420
rect 25087 3417 25099 3451
rect 25041 3411 25099 3417
rect 1452 3352 3740 3380
rect 1452 3340 1458 3352
rect 5902 3340 5908 3392
rect 5960 3340 5966 3392
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 8352 3352 8585 3380
rect 8352 3340 8358 3352
rect 8573 3349 8585 3352
rect 8619 3349 8631 3383
rect 8573 3343 8631 3349
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10413 3383 10471 3389
rect 10413 3380 10425 3383
rect 9456 3352 10425 3380
rect 9456 3340 9462 3352
rect 10413 3349 10425 3352
rect 10459 3349 10471 3383
rect 10413 3343 10471 3349
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 11977 3383 12035 3389
rect 11977 3380 11989 3383
rect 11848 3352 11989 3380
rect 11848 3340 11854 3352
rect 11977 3349 11989 3352
rect 12023 3380 12035 3383
rect 17126 3380 17132 3392
rect 12023 3352 17132 3380
rect 12023 3349 12035 3352
rect 11977 3343 12035 3349
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 21177 3383 21235 3389
rect 21177 3380 21189 3383
rect 17644 3352 21189 3380
rect 17644 3340 17650 3352
rect 21177 3349 21189 3352
rect 21223 3349 21235 3383
rect 21177 3343 21235 3349
rect 23474 3340 23480 3392
rect 23532 3380 23538 3392
rect 23845 3383 23903 3389
rect 23845 3380 23857 3383
rect 23532 3352 23857 3380
rect 23532 3340 23538 3352
rect 23845 3349 23857 3352
rect 23891 3349 23903 3383
rect 23845 3343 23903 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 1210 3136 1216 3188
rect 1268 3176 1274 3188
rect 1268 3148 2774 3176
rect 1268 3136 1274 3148
rect 1670 3068 1676 3120
rect 1728 3068 1734 3120
rect 1854 3068 1860 3120
rect 1912 3068 1918 3120
rect 2746 3108 2774 3148
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3786 3176 3792 3188
rect 3292 3148 3792 3176
rect 3292 3136 3298 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 4614 3176 4620 3188
rect 3936 3148 4620 3176
rect 3936 3136 3942 3148
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5776 3148 6193 3176
rect 5776 3136 5782 3148
rect 6181 3145 6193 3148
rect 6227 3176 6239 3179
rect 6270 3176 6276 3188
rect 6227 3148 6276 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6638 3176 6644 3188
rect 6595 3148 6644 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 6880 3148 8953 3176
rect 6880 3136 6886 3148
rect 8941 3145 8953 3148
rect 8987 3145 8999 3179
rect 8941 3139 8999 3145
rect 10042 3136 10048 3188
rect 10100 3136 10106 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 20714 3176 20720 3188
rect 18840 3148 20720 3176
rect 18840 3136 18846 3148
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 7374 3108 7380 3120
rect 2746 3080 7380 3108
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 7650 3068 7656 3120
rect 7708 3108 7714 3120
rect 8754 3108 8760 3120
rect 7708 3080 8760 3108
rect 7708 3068 7714 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 11149 3111 11207 3117
rect 11149 3108 11161 3111
rect 10008 3080 11161 3108
rect 10008 3068 10014 3080
rect 11149 3077 11161 3080
rect 11195 3077 11207 3111
rect 13372 3108 13400 3136
rect 23382 3108 23388 3120
rect 13372 3080 23388 3108
rect 11149 3071 11207 3077
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2682 3040 2688 3052
rect 2639 3012 2688 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 4890 3000 4896 3052
rect 4948 3000 4954 3052
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 6086 3040 6092 3052
rect 5215 3012 6092 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6380 3012 6745 3040
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2972 2375 2975
rect 2866 2972 2872 2984
rect 2363 2944 2872 2972
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3513 2907 3571 2913
rect 3513 2904 3525 2907
rect 2746 2876 3525 2904
rect 750 2796 756 2848
rect 808 2836 814 2848
rect 2746 2836 2774 2876
rect 3513 2873 3525 2876
rect 3559 2904 3571 2907
rect 3620 2904 3648 2935
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 6380 2981 6408 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 6972 3012 7205 3040
rect 6972 3000 6978 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 9398 3000 9404 3052
rect 9456 3000 9462 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 13173 3043 13231 3049
rect 10551 3012 13124 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 6365 2975 6423 2981
rect 6365 2972 6377 2975
rect 6236 2944 6377 2972
rect 6236 2932 6242 2944
rect 6365 2941 6377 2944
rect 6411 2941 6423 2975
rect 6365 2935 6423 2941
rect 7834 2932 7840 2984
rect 7892 2932 7898 2984
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 9950 2972 9956 2984
rect 8628 2944 9956 2972
rect 8628 2932 8634 2944
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 11698 2972 11704 2984
rect 11480 2944 11704 2972
rect 11480 2932 11486 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 10686 2904 10692 2916
rect 3559 2876 10692 2904
rect 3559 2873 3571 2876
rect 3513 2867 3571 2873
rect 10686 2864 10692 2876
rect 10744 2864 10750 2916
rect 11514 2864 11520 2916
rect 11572 2904 11578 2916
rect 11992 2904 12020 2935
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 12526 2972 12532 2984
rect 12124 2944 12532 2972
rect 12124 2932 12130 2944
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 11572 2876 12020 2904
rect 13096 2904 13124 3012
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13354 3040 13360 3052
rect 13219 3012 13360 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 16574 3040 16580 3052
rect 15059 3012 16580 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 18874 3000 18880 3052
rect 18932 3000 18938 3052
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3040 20959 3043
rect 21266 3040 21272 3052
rect 20947 3012 21272 3040
rect 20947 3009 20959 3012
rect 20901 3003 20959 3009
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 22094 3000 22100 3052
rect 22152 3000 22158 3052
rect 23842 3000 23848 3052
rect 23900 3000 23906 3052
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 16114 2904 16120 2916
rect 13096 2876 16120 2904
rect 11572 2864 11578 2876
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 19168 2904 19196 2935
rect 19518 2932 19524 2984
rect 19576 2972 19582 2984
rect 21450 2972 21456 2984
rect 19576 2944 21456 2972
rect 19576 2932 19582 2944
rect 21450 2932 21456 2944
rect 21508 2932 21514 2984
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22066 2944 22477 2972
rect 22066 2904 22094 2944
rect 22465 2941 22477 2944
rect 22511 2941 22523 2975
rect 22465 2935 22523 2941
rect 24305 2975 24363 2981
rect 24305 2941 24317 2975
rect 24351 2941 24363 2975
rect 24305 2935 24363 2941
rect 16264 2876 19196 2904
rect 19260 2876 22094 2904
rect 16264 2864 16270 2876
rect 808 2808 2774 2836
rect 808 2796 814 2808
rect 3786 2796 3792 2848
rect 3844 2836 3850 2848
rect 8294 2836 8300 2848
rect 3844 2808 8300 2836
rect 3844 2796 3850 2808
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 18230 2796 18236 2848
rect 18288 2836 18294 2848
rect 19260 2836 19288 2876
rect 18288 2808 19288 2836
rect 18288 2796 18294 2808
rect 19886 2796 19892 2848
rect 19944 2836 19950 2848
rect 24320 2836 24348 2935
rect 19944 2808 24348 2836
rect 19944 2796 19950 2808
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 1486 2592 1492 2644
rect 1544 2592 1550 2644
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 3418 2632 3424 2644
rect 2087 2604 3424 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 3568 2604 9137 2632
rect 3568 2592 3574 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13412 2604 17632 2632
rect 13412 2592 13418 2604
rect 2682 2524 2688 2576
rect 2740 2564 2746 2576
rect 4617 2567 4675 2573
rect 4617 2564 4629 2567
rect 2740 2536 4629 2564
rect 2740 2524 2746 2536
rect 4617 2533 4629 2536
rect 4663 2533 4675 2567
rect 7193 2567 7251 2573
rect 7193 2564 7205 2567
rect 4617 2527 4675 2533
rect 4816 2536 7205 2564
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 3694 2496 3700 2508
rect 2639 2468 3700 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 3344 2440 3372 2468
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 4816 2496 4844 2536
rect 7193 2533 7205 2536
rect 7239 2533 7251 2567
rect 7193 2527 7251 2533
rect 7576 2536 17540 2564
rect 3896 2468 4844 2496
rect 1946 2388 1952 2440
rect 2004 2388 2010 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 2884 2360 2912 2391
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 3896 2428 3924 2468
rect 5442 2456 5448 2508
rect 5500 2456 5506 2508
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 7576 2496 7604 2536
rect 5776 2468 7604 2496
rect 5776 2456 5782 2468
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 9030 2496 9036 2508
rect 8536 2468 9036 2496
rect 8536 2456 8542 2468
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2496 11759 2499
rect 12434 2496 12440 2508
rect 11747 2468 12440 2496
rect 11747 2465 11759 2468
rect 11701 2459 11759 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15160 2468 17325 2496
rect 15160 2456 15166 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 3660 2400 3924 2428
rect 3660 2388 3666 2400
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5810 2428 5816 2440
rect 5224 2400 5816 2428
rect 5224 2388 5230 2400
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5960 2400 6561 2428
rect 5960 2388 5966 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 7282 2360 7288 2372
rect 2884 2332 7288 2360
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7760 2304 7788 2391
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 900 2264 7665 2292
rect 900 2252 906 2264
rect 7653 2261 7665 2264
rect 7699 2292 7711 2295
rect 7742 2292 7748 2304
rect 7699 2264 7748 2292
rect 7699 2261 7711 2264
rect 7653 2255 7711 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8036 2292 8064 2391
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 17037 2431 17095 2437
rect 14691 2400 16574 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 10962 2320 10968 2372
rect 11020 2320 11026 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 15562 2360 15568 2372
rect 14016 2332 15568 2360
rect 14016 2292 14044 2332
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 16393 2363 16451 2369
rect 16393 2360 16405 2363
rect 15988 2332 16405 2360
rect 15988 2320 15994 2332
rect 16393 2329 16405 2332
rect 16439 2329 16451 2363
rect 16393 2323 16451 2329
rect 8036 2264 14044 2292
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 14918 2292 14924 2304
rect 14148 2264 14924 2292
rect 14148 2252 14154 2264
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 16080 2264 16129 2292
rect 16080 2252 16086 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16546 2292 16574 2400
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17126 2428 17132 2440
rect 17083 2400 17132 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17512 2428 17540 2536
rect 17604 2496 17632 2604
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 17736 2604 19012 2632
rect 17736 2592 17742 2604
rect 18984 2564 19012 2604
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 22278 2632 22284 2644
rect 19116 2604 22284 2632
rect 19116 2592 19122 2604
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 22370 2592 22376 2644
rect 22428 2632 22434 2644
rect 23198 2632 23204 2644
rect 22428 2604 23204 2632
rect 22428 2592 22434 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 23750 2592 23756 2644
rect 23808 2592 23814 2644
rect 24029 2635 24087 2641
rect 24029 2601 24041 2635
rect 24075 2632 24087 2635
rect 24486 2632 24492 2644
rect 24075 2604 24492 2632
rect 24075 2601 24087 2604
rect 24029 2595 24087 2601
rect 24486 2592 24492 2604
rect 24544 2592 24550 2644
rect 24578 2592 24584 2644
rect 24636 2632 24642 2644
rect 25225 2635 25283 2641
rect 25225 2632 25237 2635
rect 24636 2604 25237 2632
rect 24636 2592 24642 2604
rect 25225 2601 25237 2604
rect 25271 2601 25283 2635
rect 25225 2595 25283 2601
rect 18984 2536 22508 2564
rect 18966 2496 18972 2508
rect 17604 2468 18972 2496
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 22480 2505 22508 2536
rect 24210 2524 24216 2576
rect 24268 2524 24274 2576
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 17512 2400 18889 2428
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 19904 2360 19932 2459
rect 21453 2431 21511 2437
rect 21453 2428 21465 2431
rect 16724 2332 19932 2360
rect 21100 2400 21465 2428
rect 16724 2320 16730 2332
rect 21100 2304 21128 2400
rect 21453 2397 21465 2400
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21876 2400 22017 2428
rect 21876 2388 21882 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 18693 2295 18751 2301
rect 18693 2292 18705 2295
rect 16546 2264 18705 2292
rect 16117 2255 16175 2261
rect 18693 2261 18705 2264
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 21082 2252 21088 2304
rect 21140 2252 21146 2304
rect 21266 2252 21272 2304
rect 21324 2252 21330 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 7558 2048 7564 2100
rect 7616 2088 7622 2100
rect 8110 2088 8116 2100
rect 7616 2060 8116 2088
rect 7616 2048 7622 2060
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 11790 2020 11796 2032
rect 3476 1992 11796 2020
rect 3476 1980 3482 1992
rect 11790 1980 11796 1992
rect 11848 1980 11854 2032
rect 7190 1912 7196 1964
rect 7248 1952 7254 1964
rect 19794 1952 19800 1964
rect 7248 1924 19800 1952
rect 7248 1912 7254 1924
rect 19794 1912 19800 1924
rect 19852 1912 19858 1964
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 14090 1884 14096 1896
rect 2464 1856 14096 1884
rect 2464 1844 2470 1856
rect 14090 1844 14096 1856
rect 14148 1844 14154 1896
rect 4614 1776 4620 1828
rect 4672 1816 4678 1828
rect 10318 1816 10324 1828
rect 4672 1788 10324 1816
rect 4672 1776 4678 1788
rect 10318 1776 10324 1788
rect 10376 1776 10382 1828
rect 10962 1776 10968 1828
rect 11020 1816 11026 1828
rect 22186 1816 22192 1828
rect 11020 1788 22192 1816
rect 11020 1776 11026 1788
rect 22186 1776 22192 1788
rect 22244 1776 22250 1828
rect 5350 1708 5356 1760
rect 5408 1748 5414 1760
rect 13906 1748 13912 1760
rect 5408 1720 13912 1748
rect 5408 1708 5414 1720
rect 13906 1708 13912 1720
rect 13964 1708 13970 1760
rect 2130 1640 2136 1692
rect 2188 1680 2194 1692
rect 17494 1680 17500 1692
rect 2188 1652 17500 1680
rect 2188 1640 2194 1652
rect 17494 1640 17500 1652
rect 17552 1640 17558 1692
rect 5258 1572 5264 1624
rect 5316 1612 5322 1624
rect 9766 1612 9772 1624
rect 5316 1584 9772 1612
rect 5316 1572 5322 1584
rect 9766 1572 9772 1584
rect 9824 1572 9830 1624
rect 9490 1504 9496 1556
rect 9548 1544 9554 1556
rect 24578 1544 24584 1556
rect 9548 1516 24584 1544
rect 9548 1504 9554 1516
rect 24578 1504 24584 1516
rect 24636 1504 24642 1556
rect 9306 1436 9312 1488
rect 9364 1476 9370 1488
rect 17218 1476 17224 1488
rect 9364 1448 17224 1476
rect 9364 1436 9370 1448
rect 17218 1436 17224 1448
rect 17276 1436 17282 1488
rect 1762 1368 1768 1420
rect 1820 1408 1826 1420
rect 9582 1408 9588 1420
rect 1820 1380 9588 1408
rect 1820 1368 1826 1380
rect 9582 1368 9588 1380
rect 9640 1368 9646 1420
rect 7926 1300 7932 1352
rect 7984 1340 7990 1352
rect 24394 1340 24400 1352
rect 7984 1312 24400 1340
rect 7984 1300 7990 1312
rect 24394 1300 24400 1312
rect 24452 1300 24458 1352
rect 8662 1232 8668 1284
rect 8720 1272 8726 1284
rect 21266 1272 21272 1284
rect 8720 1244 21272 1272
rect 8720 1232 8726 1244
rect 21266 1232 21272 1244
rect 21324 1232 21330 1284
rect 6454 1164 6460 1216
rect 6512 1204 6518 1216
rect 20070 1204 20076 1216
rect 6512 1176 20076 1204
rect 6512 1164 6518 1176
rect 20070 1164 20076 1176
rect 20128 1164 20134 1216
rect 4154 1096 4160 1148
rect 4212 1136 4218 1148
rect 18874 1136 18880 1148
rect 4212 1108 18880 1136
rect 4212 1096 4218 1108
rect 18874 1096 18880 1108
rect 18932 1096 18938 1148
rect 8294 1028 8300 1080
rect 8352 1068 8358 1080
rect 21082 1068 21088 1080
rect 8352 1040 21088 1068
rect 8352 1028 8358 1040
rect 21082 1028 21088 1040
rect 21140 1028 21146 1080
rect 7834 960 7840 1012
rect 7892 1000 7898 1012
rect 19610 1000 19616 1012
rect 7892 972 19616 1000
rect 7892 960 7898 972
rect 19610 960 19616 972
rect 19668 960 19674 1012
rect 7650 892 7656 944
rect 7708 932 7714 944
rect 20898 932 20904 944
rect 7708 904 20904 932
rect 7708 892 7714 904
rect 20898 892 20904 904
rect 20956 892 20962 944
rect 7466 824 7472 876
rect 7524 864 7530 876
rect 19702 864 19708 876
rect 7524 836 19708 864
rect 7524 824 7530 836
rect 19702 824 19708 836
rect 19760 824 19766 876
rect 4338 144 4344 196
rect 4396 184 4402 196
rect 12434 184 12440 196
rect 4396 156 12440 184
rect 4396 144 4402 156
rect 12434 144 12440 156
rect 12492 144 12498 196
rect 6178 76 6184 128
rect 6236 116 6242 128
rect 24210 116 24216 128
rect 6236 88 24216 116
rect 6236 76 6242 88
rect 24210 76 24216 88
rect 24268 76 24274 128
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 18972 54315 19024 54324
rect 18972 54281 18981 54315
rect 18981 54281 19015 54315
rect 19015 54281 19024 54315
rect 18972 54272 19024 54281
rect 3884 54136 3936 54188
rect 6552 54136 6604 54188
rect 6736 54179 6788 54188
rect 6736 54145 6745 54179
rect 6745 54145 6779 54179
rect 6779 54145 6788 54179
rect 6736 54136 6788 54145
rect 13452 54136 13504 54188
rect 14832 54136 14884 54188
rect 16580 54136 16632 54188
rect 17592 54136 17644 54188
rect 25320 54204 25372 54256
rect 2412 54068 2464 54120
rect 4068 54068 4120 54120
rect 6920 54068 6972 54120
rect 11060 54068 11112 54120
rect 18972 54068 19024 54120
rect 16764 54000 16816 54052
rect 25228 54136 25280 54188
rect 25136 54068 25188 54120
rect 23388 54000 23440 54052
rect 23480 54000 23532 54052
rect 13544 53975 13596 53984
rect 13544 53941 13553 53975
rect 13553 53941 13587 53975
rect 13587 53941 13596 53975
rect 13544 53932 13596 53941
rect 14924 53975 14976 53984
rect 14924 53941 14933 53975
rect 14933 53941 14967 53975
rect 14967 53941 14976 53975
rect 14924 53932 14976 53941
rect 15660 53932 15712 53984
rect 17132 53932 17184 53984
rect 23940 53932 23992 53984
rect 24584 53932 24636 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 25228 53771 25280 53780
rect 25228 53737 25237 53771
rect 25237 53737 25271 53771
rect 25271 53737 25280 53771
rect 25228 53728 25280 53737
rect 24860 53660 24912 53712
rect 25872 53660 25924 53712
rect 1032 53592 1084 53644
rect 5172 53592 5224 53644
rect 7656 53524 7708 53576
rect 22376 53567 22428 53576
rect 22376 53533 22385 53567
rect 22385 53533 22419 53567
rect 22419 53533 22428 53567
rect 22376 53524 22428 53533
rect 23296 53524 23348 53576
rect 24584 53567 24636 53576
rect 24584 53533 24593 53567
rect 24593 53533 24627 53567
rect 24627 53533 24636 53567
rect 24584 53524 24636 53533
rect 5540 53456 5592 53508
rect 22100 53388 22152 53440
rect 23756 53431 23808 53440
rect 23756 53397 23765 53431
rect 23765 53397 23799 53431
rect 23799 53397 23808 53431
rect 23756 53388 23808 53397
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 3884 53184 3936 53236
rect 6552 53227 6604 53236
rect 6552 53193 6561 53227
rect 6561 53193 6595 53227
rect 6595 53193 6604 53227
rect 6552 53184 6604 53193
rect 25136 53184 25188 53236
rect 22836 53159 22888 53168
rect 22836 53125 22845 53159
rect 22845 53125 22879 53159
rect 22879 53125 22888 53159
rect 22836 53116 22888 53125
rect 8852 53048 8904 53100
rect 16212 53048 16264 53100
rect 20352 53048 20404 53100
rect 24860 53116 24912 53168
rect 23940 53048 23992 53100
rect 7748 52980 7800 53032
rect 18972 52912 19024 52964
rect 24676 52844 24728 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 7656 52683 7708 52692
rect 7656 52649 7665 52683
rect 7665 52649 7699 52683
rect 7699 52649 7708 52683
rect 7656 52640 7708 52649
rect 23296 52640 23348 52692
rect 25320 52683 25372 52692
rect 25320 52649 25329 52683
rect 25329 52649 25363 52683
rect 25363 52649 25372 52683
rect 25320 52640 25372 52649
rect 7840 52572 7892 52624
rect 8392 52572 8444 52624
rect 9588 52436 9640 52488
rect 17224 52436 17276 52488
rect 22744 52436 22796 52488
rect 23480 52436 23532 52488
rect 24124 52436 24176 52488
rect 24676 52479 24728 52488
rect 24676 52445 24685 52479
rect 24685 52445 24719 52479
rect 24719 52445 24728 52479
rect 24676 52436 24728 52445
rect 23940 52343 23992 52352
rect 23940 52309 23949 52343
rect 23949 52309 23983 52343
rect 23983 52309 23992 52343
rect 23940 52300 23992 52309
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 6736 52096 6788 52148
rect 24952 52071 25004 52080
rect 24952 52037 24961 52071
rect 24961 52037 24995 52071
rect 24995 52037 25004 52071
rect 24952 52028 25004 52037
rect 10784 51960 10836 52012
rect 23756 51960 23808 52012
rect 24584 51960 24636 52012
rect 18696 51892 18748 51944
rect 17316 51824 17368 51876
rect 22560 51756 22612 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 24124 51595 24176 51604
rect 24124 51561 24133 51595
rect 24133 51561 24167 51595
rect 24167 51561 24176 51595
rect 24124 51552 24176 51561
rect 24584 51595 24636 51604
rect 24584 51561 24593 51595
rect 24593 51561 24627 51595
rect 24627 51561 24636 51595
rect 24584 51552 24636 51561
rect 24952 51484 25004 51536
rect 24952 51323 25004 51332
rect 24952 51289 24961 51323
rect 24961 51289 24995 51323
rect 24995 51289 25004 51323
rect 24952 51280 25004 51289
rect 25044 51255 25096 51264
rect 25044 51221 25053 51255
rect 25053 51221 25087 51255
rect 25087 51221 25096 51255
rect 25044 51212 25096 51221
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 7748 51008 7800 51060
rect 5540 50668 5592 50720
rect 6828 50668 6880 50720
rect 24952 50915 25004 50924
rect 24952 50881 24961 50915
rect 24961 50881 24995 50915
rect 24995 50881 25004 50915
rect 24952 50872 25004 50881
rect 11060 50668 11112 50720
rect 24584 50668 24636 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 16396 50464 16448 50516
rect 24584 50464 24636 50516
rect 6828 50328 6880 50380
rect 8300 50328 8352 50380
rect 16488 50328 16540 50380
rect 24492 50328 24544 50380
rect 25504 50167 25556 50176
rect 25504 50133 25513 50167
rect 25513 50133 25547 50167
rect 25547 50133 25556 50167
rect 25504 50124 25556 50133
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 25504 49784 25556 49836
rect 24768 49759 24820 49768
rect 24768 49725 24777 49759
rect 24777 49725 24811 49759
rect 24811 49725 24820 49759
rect 24768 49716 24820 49725
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 18788 49376 18840 49428
rect 22100 49376 22152 49428
rect 22560 49215 22612 49224
rect 22560 49181 22569 49215
rect 22569 49181 22603 49215
rect 22603 49181 22612 49215
rect 22560 49172 22612 49181
rect 25136 49147 25188 49156
rect 25136 49113 25145 49147
rect 25145 49113 25179 49147
rect 25179 49113 25188 49147
rect 25136 49104 25188 49113
rect 22652 49036 22704 49088
rect 25228 49079 25280 49088
rect 25228 49045 25237 49079
rect 25237 49045 25271 49079
rect 25271 49045 25280 49079
rect 25228 49036 25280 49045
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 8852 48832 8904 48884
rect 11428 48832 11480 48884
rect 7748 48764 7800 48816
rect 8208 48764 8260 48816
rect 11060 48764 11112 48816
rect 7748 48671 7800 48680
rect 7748 48637 7757 48671
rect 7757 48637 7791 48671
rect 7791 48637 7800 48671
rect 7748 48628 7800 48637
rect 8392 48671 8444 48680
rect 8392 48637 8401 48671
rect 8401 48637 8435 48671
rect 8435 48637 8444 48671
rect 8392 48628 8444 48637
rect 10140 48535 10192 48544
rect 10140 48501 10149 48535
rect 10149 48501 10183 48535
rect 10183 48501 10192 48535
rect 10140 48492 10192 48501
rect 25136 48492 25188 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 8300 48263 8352 48272
rect 8300 48229 8309 48263
rect 8309 48229 8343 48263
rect 8343 48229 8352 48263
rect 8300 48220 8352 48229
rect 8576 48152 8628 48204
rect 8208 48084 8260 48136
rect 9128 48127 9180 48136
rect 9128 48093 9137 48127
rect 9137 48093 9171 48127
rect 9171 48093 9180 48127
rect 9128 48084 9180 48093
rect 11428 48127 11480 48136
rect 11428 48093 11472 48127
rect 11472 48093 11480 48127
rect 11428 48084 11480 48093
rect 25136 48127 25188 48136
rect 25136 48093 25145 48127
rect 25145 48093 25179 48127
rect 25179 48093 25188 48127
rect 25136 48084 25188 48093
rect 7840 48016 7892 48068
rect 8576 47991 8628 48000
rect 8576 47957 8585 47991
rect 8585 47957 8619 47991
rect 8619 47957 8628 47991
rect 8576 47948 8628 47957
rect 11428 47948 11480 48000
rect 14464 47948 14516 48000
rect 24860 47948 24912 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 8852 47719 8904 47728
rect 8852 47685 8861 47719
rect 8861 47685 8895 47719
rect 8895 47685 8904 47719
rect 8852 47676 8904 47685
rect 9312 47583 9364 47592
rect 9312 47549 9321 47583
rect 9321 47549 9355 47583
rect 9355 47549 9364 47583
rect 9312 47540 9364 47549
rect 9588 47540 9640 47592
rect 25320 47651 25372 47660
rect 25320 47617 25329 47651
rect 25329 47617 25363 47651
rect 25363 47617 25372 47651
rect 25320 47608 25372 47617
rect 8760 47472 8812 47524
rect 7840 47404 7892 47456
rect 10508 47404 10560 47456
rect 14648 47404 14700 47456
rect 25780 47404 25832 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 9128 47200 9180 47252
rect 10324 47243 10376 47252
rect 10324 47209 10333 47243
rect 10333 47209 10367 47243
rect 10367 47209 10376 47243
rect 10324 47200 10376 47209
rect 11060 47243 11112 47252
rect 11060 47209 11069 47243
rect 11069 47209 11103 47243
rect 11103 47209 11112 47243
rect 11060 47200 11112 47209
rect 9588 47132 9640 47184
rect 14924 47064 14976 47116
rect 9772 46996 9824 47048
rect 11060 46996 11112 47048
rect 12164 46996 12216 47048
rect 22652 47039 22704 47048
rect 22652 47005 22661 47039
rect 22661 47005 22695 47039
rect 22695 47005 22704 47039
rect 22652 46996 22704 47005
rect 14280 46928 14332 46980
rect 14464 46971 14516 46980
rect 14464 46937 14473 46971
rect 14473 46937 14507 46971
rect 14507 46937 14516 46971
rect 14464 46928 14516 46937
rect 20444 46928 20496 46980
rect 20812 46928 20864 46980
rect 25320 46860 25372 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 11428 46588 11480 46640
rect 14648 46631 14700 46640
rect 14648 46597 14657 46631
rect 14657 46597 14691 46631
rect 14691 46597 14700 46631
rect 14648 46588 14700 46597
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 13544 46452 13596 46504
rect 15660 46452 15712 46504
rect 21732 46452 21784 46504
rect 19708 46384 19760 46436
rect 22652 46316 22704 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 9772 46155 9824 46164
rect 9772 46121 9781 46155
rect 9781 46121 9815 46155
rect 9815 46121 9824 46155
rect 9772 46112 9824 46121
rect 10140 45976 10192 46028
rect 10784 46019 10836 46028
rect 10784 45985 10793 46019
rect 10793 45985 10827 46019
rect 10827 45985 10836 46019
rect 10784 45976 10836 45985
rect 12072 46019 12124 46028
rect 12072 45985 12081 46019
rect 12081 45985 12115 46019
rect 12115 45985 12124 46019
rect 12072 45976 12124 45985
rect 14280 45976 14332 46028
rect 9312 45908 9364 45960
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 17132 45840 17184 45892
rect 20168 45840 20220 45892
rect 22468 45772 22520 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 10784 45568 10836 45620
rect 12164 45611 12216 45620
rect 12164 45577 12173 45611
rect 12173 45577 12207 45611
rect 12207 45577 12216 45611
rect 12164 45568 12216 45577
rect 9496 45543 9548 45552
rect 9496 45509 9505 45543
rect 9505 45509 9539 45543
rect 9539 45509 9548 45543
rect 9496 45500 9548 45509
rect 11152 45432 11204 45484
rect 9036 45364 9088 45416
rect 10968 45407 11020 45416
rect 10968 45373 10977 45407
rect 10977 45373 11011 45407
rect 11011 45373 11020 45407
rect 10968 45364 11020 45373
rect 11796 45271 11848 45280
rect 11796 45237 11805 45271
rect 11805 45237 11839 45271
rect 11839 45237 11848 45271
rect 11796 45228 11848 45237
rect 25320 45228 25372 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 10140 45024 10192 45076
rect 8576 44888 8628 44940
rect 11520 44888 11572 44940
rect 10508 44820 10560 44872
rect 10876 44820 10928 44872
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 22376 44684 22428 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 10876 44523 10928 44532
rect 10876 44489 10885 44523
rect 10885 44489 10919 44523
rect 10919 44489 10928 44523
rect 10876 44480 10928 44489
rect 10232 44387 10284 44396
rect 10232 44353 10241 44387
rect 10241 44353 10275 44387
rect 10275 44353 10284 44387
rect 10232 44344 10284 44353
rect 24768 44387 24820 44396
rect 24768 44353 24777 44387
rect 24777 44353 24811 44387
rect 24811 44353 24820 44387
rect 24768 44344 24820 44353
rect 11520 44276 11572 44328
rect 14372 44208 14424 44260
rect 10508 44140 10560 44192
rect 11980 44140 12032 44192
rect 19064 44140 19116 44192
rect 25044 44140 25096 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 10232 43936 10284 43988
rect 20812 43843 20864 43852
rect 20812 43809 20821 43843
rect 20821 43809 20855 43843
rect 20855 43809 20864 43843
rect 20812 43800 20864 43809
rect 21272 43800 21324 43852
rect 9956 43775 10008 43784
rect 9956 43741 9965 43775
rect 9965 43741 9999 43775
rect 9999 43741 10008 43775
rect 9956 43732 10008 43741
rect 10324 43732 10376 43784
rect 19432 43732 19484 43784
rect 11980 43664 12032 43716
rect 21088 43664 21140 43716
rect 21272 43664 21324 43716
rect 20628 43596 20680 43648
rect 25504 43639 25556 43648
rect 25504 43605 25513 43639
rect 25513 43605 25547 43639
rect 25547 43605 25556 43639
rect 25504 43596 25556 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 25504 43324 25556 43376
rect 23480 43052 23532 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 11888 42848 11940 42900
rect 11520 42712 11572 42764
rect 11980 42755 12032 42764
rect 11980 42721 11989 42755
rect 11989 42721 12023 42755
rect 12023 42721 12032 42755
rect 11980 42712 12032 42721
rect 15936 42712 15988 42764
rect 17316 42712 17368 42764
rect 25136 42619 25188 42628
rect 25136 42585 25145 42619
rect 25145 42585 25179 42619
rect 25179 42585 25188 42619
rect 25136 42576 25188 42585
rect 9956 42508 10008 42560
rect 11520 42508 11572 42560
rect 25228 42551 25280 42560
rect 25228 42517 25237 42551
rect 25237 42517 25271 42551
rect 25271 42517 25280 42551
rect 25228 42508 25280 42517
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 25320 41964 25372 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 25136 41531 25188 41540
rect 25136 41497 25145 41531
rect 25145 41497 25179 41531
rect 25179 41497 25188 41531
rect 25136 41488 25188 41497
rect 16672 41420 16724 41472
rect 23940 41420 23992 41472
rect 24860 41420 24912 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 17224 41080 17276 41132
rect 20628 41080 20680 41132
rect 24860 41080 24912 41132
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 18328 40876 18380 40928
rect 23848 40876 23900 40928
rect 24952 40876 25004 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 24676 40375 24728 40384
rect 24676 40341 24685 40375
rect 24685 40341 24719 40375
rect 24719 40341 24728 40375
rect 24676 40332 24728 40341
rect 24768 40332 24820 40384
rect 26148 40332 26200 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 24768 40060 24820 40112
rect 24860 39992 24912 40044
rect 17040 39856 17092 39908
rect 24400 39831 24452 39840
rect 24400 39797 24409 39831
rect 24409 39797 24443 39831
rect 24443 39797 24452 39831
rect 24400 39788 24452 39797
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 11888 39627 11940 39636
rect 11888 39593 11897 39627
rect 11897 39593 11931 39627
rect 11931 39593 11940 39627
rect 11888 39584 11940 39593
rect 24860 39584 24912 39636
rect 11244 39423 11296 39432
rect 11244 39389 11253 39423
rect 11253 39389 11287 39423
rect 11287 39389 11296 39423
rect 11244 39380 11296 39389
rect 24308 39312 24360 39364
rect 25504 39312 25556 39364
rect 24492 39287 24544 39296
rect 24492 39253 24501 39287
rect 24501 39253 24535 39287
rect 24535 39253 24544 39287
rect 24492 39244 24544 39253
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 7748 39040 7800 39092
rect 8852 38904 8904 38956
rect 24492 38904 24544 38956
rect 25136 38904 25188 38956
rect 21088 38700 21140 38752
rect 25320 38743 25372 38752
rect 25320 38709 25329 38743
rect 25329 38709 25363 38743
rect 25363 38709 25372 38743
rect 25320 38700 25372 38709
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 20076 38428 20128 38480
rect 18328 38292 18380 38344
rect 14556 38156 14608 38208
rect 22744 38156 22796 38208
rect 24584 38335 24636 38344
rect 24584 38301 24593 38335
rect 24593 38301 24627 38335
rect 24627 38301 24636 38335
rect 24584 38292 24636 38301
rect 24952 38156 25004 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 11244 37952 11296 38004
rect 11152 37816 11204 37868
rect 11796 37816 11848 37868
rect 17316 37816 17368 37868
rect 23664 37816 23716 37868
rect 25044 37680 25096 37732
rect 23480 37612 23532 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 23480 37204 23532 37256
rect 25228 37204 25280 37256
rect 22192 37068 22244 37120
rect 25412 37068 25464 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 20444 36864 20496 36916
rect 24584 36864 24636 36916
rect 22284 36771 22336 36780
rect 22284 36737 22293 36771
rect 22293 36737 22327 36771
rect 22327 36737 22336 36771
rect 22284 36728 22336 36737
rect 25320 36796 25372 36848
rect 24768 36728 24820 36780
rect 23388 36524 23440 36576
rect 24584 36524 24636 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 22284 36320 22336 36372
rect 25228 36363 25280 36372
rect 25228 36329 25237 36363
rect 25237 36329 25271 36363
rect 25271 36329 25280 36363
rect 25228 36320 25280 36329
rect 19984 36159 20036 36168
rect 19984 36125 19993 36159
rect 19993 36125 20027 36159
rect 20027 36125 20036 36159
rect 19984 36116 20036 36125
rect 21456 36116 21508 36168
rect 23296 36159 23348 36168
rect 23296 36125 23305 36159
rect 23305 36125 23339 36159
rect 23339 36125 23348 36159
rect 23296 36116 23348 36125
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 24216 36048 24268 36100
rect 23204 35980 23256 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 8760 35819 8812 35828
rect 8760 35785 8769 35819
rect 8769 35785 8803 35819
rect 8803 35785 8812 35819
rect 8760 35776 8812 35785
rect 9128 35640 9180 35692
rect 11520 35776 11572 35828
rect 20444 35776 20496 35828
rect 11704 35751 11756 35760
rect 11704 35717 11713 35751
rect 11713 35717 11747 35751
rect 11747 35717 11756 35751
rect 11704 35708 11756 35717
rect 19156 35640 19208 35692
rect 22468 35819 22520 35828
rect 22468 35785 22477 35819
rect 22477 35785 22511 35819
rect 22511 35785 22520 35819
rect 22468 35776 22520 35785
rect 22652 35708 22704 35760
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 11152 35615 11204 35624
rect 11152 35581 11161 35615
rect 11161 35581 11195 35615
rect 11195 35581 11204 35615
rect 11152 35572 11204 35581
rect 21180 35572 21232 35624
rect 21732 35640 21784 35692
rect 22560 35615 22612 35624
rect 22560 35581 22569 35615
rect 22569 35581 22603 35615
rect 22603 35581 22612 35615
rect 22560 35572 22612 35581
rect 23204 35683 23256 35692
rect 23204 35649 23213 35683
rect 23213 35649 23247 35683
rect 23247 35649 23256 35683
rect 23204 35640 23256 35649
rect 23388 35640 23440 35692
rect 25872 35572 25924 35624
rect 20812 35504 20864 35556
rect 11612 35479 11664 35488
rect 11612 35445 11621 35479
rect 11621 35445 11655 35479
rect 11655 35445 11664 35479
rect 11612 35436 11664 35445
rect 20260 35479 20312 35488
rect 20260 35445 20269 35479
rect 20269 35445 20303 35479
rect 20303 35445 20312 35479
rect 20260 35436 20312 35445
rect 20720 35479 20772 35488
rect 20720 35445 20729 35479
rect 20729 35445 20763 35479
rect 20763 35445 20772 35479
rect 20720 35436 20772 35445
rect 20996 35436 21048 35488
rect 23940 35436 23992 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 22284 35232 22336 35284
rect 21732 35207 21784 35216
rect 21732 35173 21741 35207
rect 21741 35173 21775 35207
rect 21775 35173 21784 35207
rect 21732 35164 21784 35173
rect 22652 35164 22704 35216
rect 20168 35096 20220 35148
rect 19524 35028 19576 35080
rect 20260 35028 20312 35080
rect 21824 34960 21876 35012
rect 22376 35096 22428 35148
rect 23296 35139 23348 35148
rect 23296 35105 23305 35139
rect 23305 35105 23339 35139
rect 23339 35105 23348 35139
rect 23296 35096 23348 35105
rect 23388 35028 23440 35080
rect 25228 35028 25280 35080
rect 24308 34960 24360 35012
rect 18328 34892 18380 34944
rect 19616 34892 19668 34944
rect 20352 34892 20404 34944
rect 22468 34892 22520 34944
rect 23388 34892 23440 34944
rect 24032 34892 24084 34944
rect 24952 34892 25004 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 19156 34731 19208 34740
rect 19156 34697 19165 34731
rect 19165 34697 19199 34731
rect 19199 34697 19208 34731
rect 19156 34688 19208 34697
rect 19708 34688 19760 34740
rect 21180 34620 21232 34672
rect 19616 34595 19668 34604
rect 19616 34561 19625 34595
rect 19625 34561 19659 34595
rect 19659 34561 19668 34595
rect 19616 34552 19668 34561
rect 21364 34552 21416 34604
rect 22836 34552 22888 34604
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 18328 34484 18380 34536
rect 17040 34416 17092 34468
rect 22652 34527 22704 34536
rect 22652 34493 22661 34527
rect 22661 34493 22695 34527
rect 22695 34493 22704 34527
rect 22652 34484 22704 34493
rect 23756 34527 23808 34536
rect 23756 34493 23765 34527
rect 23765 34493 23799 34527
rect 23799 34493 23808 34527
rect 23756 34484 23808 34493
rect 24860 34484 24912 34536
rect 25320 34484 25372 34536
rect 19892 34348 19944 34400
rect 22100 34416 22152 34468
rect 22560 34416 22612 34468
rect 23388 34348 23440 34400
rect 24860 34391 24912 34400
rect 24860 34357 24869 34391
rect 24869 34357 24903 34391
rect 24903 34357 24912 34391
rect 24860 34348 24912 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 9680 34144 9732 34196
rect 24860 34144 24912 34196
rect 25228 34187 25280 34196
rect 25228 34153 25237 34187
rect 25237 34153 25271 34187
rect 25271 34153 25280 34187
rect 25228 34144 25280 34153
rect 21180 34119 21232 34128
rect 21180 34085 21189 34119
rect 21189 34085 21223 34119
rect 21223 34085 21232 34119
rect 21180 34076 21232 34085
rect 23388 34119 23440 34128
rect 23388 34085 23397 34119
rect 23397 34085 23431 34119
rect 23431 34085 23440 34119
rect 23388 34076 23440 34085
rect 11612 34008 11664 34060
rect 19432 34051 19484 34060
rect 19432 34017 19441 34051
rect 19441 34017 19475 34051
rect 19475 34017 19484 34051
rect 21640 34051 21692 34060
rect 19432 34008 19484 34017
rect 21640 34017 21649 34051
rect 21649 34017 21683 34051
rect 21683 34017 21692 34051
rect 21640 34008 21692 34017
rect 9772 33983 9824 33992
rect 9772 33949 9781 33983
rect 9781 33949 9815 33983
rect 9815 33949 9824 33983
rect 9772 33940 9824 33949
rect 17040 33983 17092 33992
rect 17040 33949 17049 33983
rect 17049 33949 17083 33983
rect 17083 33949 17092 33983
rect 17040 33940 17092 33949
rect 18328 33940 18380 33992
rect 24032 33983 24084 33992
rect 24032 33949 24041 33983
rect 24041 33949 24075 33983
rect 24075 33949 24084 33983
rect 24032 33940 24084 33949
rect 25688 33940 25740 33992
rect 15384 33872 15436 33924
rect 18512 33804 18564 33856
rect 21180 33872 21232 33924
rect 22192 33872 22244 33924
rect 21456 33804 21508 33856
rect 22008 33804 22060 33856
rect 25596 33804 25648 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 16212 33643 16264 33652
rect 16212 33609 16221 33643
rect 16221 33609 16255 33643
rect 16255 33609 16264 33643
rect 16212 33600 16264 33609
rect 16488 33643 16540 33652
rect 16488 33609 16497 33643
rect 16497 33609 16531 33643
rect 16531 33609 16540 33643
rect 16488 33600 16540 33609
rect 18328 33600 18380 33652
rect 19984 33600 20036 33652
rect 20444 33600 20496 33652
rect 18420 33464 18472 33516
rect 19340 33464 19392 33516
rect 20904 33464 20956 33516
rect 21180 33464 21232 33516
rect 22008 33600 22060 33652
rect 21640 33532 21692 33584
rect 22284 33532 22336 33584
rect 23848 33600 23900 33652
rect 25228 33600 25280 33652
rect 25872 33600 25924 33652
rect 24584 33507 24636 33516
rect 24584 33473 24593 33507
rect 24593 33473 24627 33507
rect 24627 33473 24636 33507
rect 24584 33464 24636 33473
rect 19432 33396 19484 33448
rect 20812 33396 20864 33448
rect 23940 33396 23992 33448
rect 24768 33439 24820 33448
rect 24768 33405 24777 33439
rect 24777 33405 24811 33439
rect 24811 33405 24820 33439
rect 24768 33396 24820 33405
rect 19248 33260 19300 33312
rect 22008 33260 22060 33312
rect 23480 33260 23532 33312
rect 23664 33260 23716 33312
rect 24216 33303 24268 33312
rect 24216 33269 24225 33303
rect 24225 33269 24259 33303
rect 24259 33269 24268 33303
rect 24216 33260 24268 33269
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 9312 33099 9364 33108
rect 9312 33065 9321 33099
rect 9321 33065 9355 33099
rect 9355 33065 9364 33099
rect 9312 33056 9364 33065
rect 18420 33099 18472 33108
rect 18420 33065 18429 33099
rect 18429 33065 18463 33099
rect 18463 33065 18472 33099
rect 18420 33056 18472 33065
rect 18696 33099 18748 33108
rect 18696 33065 18705 33099
rect 18705 33065 18739 33099
rect 18739 33065 18748 33099
rect 18696 33056 18748 33065
rect 18972 33099 19024 33108
rect 18972 33065 18981 33099
rect 18981 33065 19015 33099
rect 19015 33065 19024 33099
rect 18972 33056 19024 33065
rect 19340 33056 19392 33108
rect 22100 33056 22152 33108
rect 23204 33056 23256 33108
rect 23296 33056 23348 33108
rect 17224 32963 17276 32972
rect 17224 32929 17233 32963
rect 17233 32929 17267 32963
rect 17267 32929 17276 32963
rect 17224 32920 17276 32929
rect 20904 32988 20956 33040
rect 21364 32988 21416 33040
rect 7748 32852 7800 32904
rect 16488 32852 16540 32904
rect 17592 32852 17644 32904
rect 20352 32920 20404 32972
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 22928 32920 22980 32972
rect 24400 32920 24452 32972
rect 18788 32852 18840 32904
rect 19432 32895 19484 32904
rect 19432 32861 19441 32895
rect 19441 32861 19475 32895
rect 19475 32861 19484 32895
rect 19432 32852 19484 32861
rect 20812 32852 20864 32904
rect 16212 32784 16264 32836
rect 16856 32784 16908 32836
rect 18604 32784 18656 32836
rect 14740 32716 14792 32768
rect 16580 32759 16632 32768
rect 16580 32725 16589 32759
rect 16589 32725 16623 32759
rect 16623 32725 16632 32759
rect 16580 32716 16632 32725
rect 18420 32716 18472 32768
rect 22008 32852 22060 32904
rect 25228 32852 25280 32904
rect 23020 32784 23072 32836
rect 21640 32759 21692 32768
rect 21640 32725 21649 32759
rect 21649 32725 21683 32759
rect 21683 32725 21692 32759
rect 21640 32716 21692 32725
rect 23204 32716 23256 32768
rect 25044 32784 25096 32836
rect 23940 32716 23992 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 9036 32555 9088 32564
rect 9036 32521 9045 32555
rect 9045 32521 9079 32555
rect 9079 32521 9088 32555
rect 9036 32512 9088 32521
rect 15384 32487 15436 32496
rect 15384 32453 15393 32487
rect 15393 32453 15427 32487
rect 15427 32453 15436 32487
rect 15384 32444 15436 32453
rect 18420 32444 18472 32496
rect 25044 32512 25096 32564
rect 21456 32444 21508 32496
rect 22284 32444 22336 32496
rect 9220 32419 9272 32428
rect 9220 32385 9229 32419
rect 9229 32385 9263 32419
rect 9263 32385 9272 32419
rect 9220 32376 9272 32385
rect 23020 32444 23072 32496
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 14280 32308 14332 32360
rect 17132 32308 17184 32360
rect 18512 32308 18564 32360
rect 19432 32308 19484 32360
rect 20628 32351 20680 32360
rect 20628 32317 20637 32351
rect 20637 32317 20671 32351
rect 20671 32317 20680 32351
rect 20628 32308 20680 32317
rect 25412 32308 25464 32360
rect 15016 32172 15068 32224
rect 19524 32172 19576 32224
rect 22560 32172 22612 32224
rect 25136 32215 25188 32224
rect 25136 32181 25145 32215
rect 25145 32181 25179 32215
rect 25179 32181 25188 32215
rect 25136 32172 25188 32181
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 9772 31968 9824 32020
rect 13912 31968 13964 32020
rect 16672 32011 16724 32020
rect 16672 31977 16681 32011
rect 16681 31977 16715 32011
rect 16715 31977 16724 32011
rect 16672 31968 16724 31977
rect 12072 31900 12124 31952
rect 16948 31900 17000 31952
rect 10508 31832 10560 31884
rect 12624 31832 12676 31884
rect 14280 31875 14332 31884
rect 14280 31841 14289 31875
rect 14289 31841 14323 31875
rect 14323 31841 14332 31875
rect 14280 31832 14332 31841
rect 14556 31875 14608 31884
rect 14556 31841 14565 31875
rect 14565 31841 14599 31875
rect 14599 31841 14608 31875
rect 14556 31832 14608 31841
rect 19432 31968 19484 32020
rect 20812 31968 20864 32020
rect 21456 32011 21508 32020
rect 21456 31977 21465 32011
rect 21465 31977 21499 32011
rect 21499 31977 21508 32011
rect 21456 31968 21508 31977
rect 21640 31968 21692 32020
rect 25412 31968 25464 32020
rect 18788 31943 18840 31952
rect 18788 31909 18797 31943
rect 18797 31909 18831 31943
rect 18831 31909 18840 31943
rect 18788 31900 18840 31909
rect 24860 31900 24912 31952
rect 9680 31764 9732 31816
rect 11152 31764 11204 31816
rect 14004 31764 14056 31816
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 13544 31696 13596 31748
rect 15016 31696 15068 31748
rect 18696 31696 18748 31748
rect 19708 31739 19760 31748
rect 19708 31705 19717 31739
rect 19717 31705 19751 31739
rect 19751 31705 19760 31739
rect 19708 31696 19760 31705
rect 20536 31628 20588 31680
rect 21640 31807 21692 31816
rect 21640 31773 21649 31807
rect 21649 31773 21683 31807
rect 21683 31773 21692 31807
rect 21640 31764 21692 31773
rect 21824 31832 21876 31884
rect 22560 31875 22612 31884
rect 22560 31841 22569 31875
rect 22569 31841 22603 31875
rect 22603 31841 22612 31875
rect 22560 31832 22612 31841
rect 25320 31832 25372 31884
rect 23204 31807 23256 31816
rect 23204 31773 23213 31807
rect 23213 31773 23247 31807
rect 23247 31773 23256 31807
rect 23204 31764 23256 31773
rect 25228 31764 25280 31816
rect 24768 31628 24820 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 19708 31424 19760 31476
rect 20168 31424 20220 31476
rect 20260 31424 20312 31476
rect 21456 31424 21508 31476
rect 23204 31424 23256 31476
rect 24676 31424 24728 31476
rect 11244 31288 11296 31340
rect 13912 31288 13964 31340
rect 14556 31331 14608 31340
rect 14556 31297 14565 31331
rect 14565 31297 14599 31331
rect 14599 31297 14608 31331
rect 14556 31288 14608 31297
rect 23940 31356 23992 31408
rect 24124 31356 24176 31408
rect 17868 31288 17920 31340
rect 19616 31263 19668 31272
rect 19616 31229 19625 31263
rect 19625 31229 19659 31263
rect 19659 31229 19668 31263
rect 19616 31220 19668 31229
rect 19708 31220 19760 31272
rect 22008 31331 22060 31340
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 23388 31331 23440 31340
rect 23388 31297 23397 31331
rect 23397 31297 23431 31331
rect 23431 31297 23440 31331
rect 23388 31288 23440 31297
rect 10324 31152 10376 31204
rect 21364 31152 21416 31204
rect 9772 31084 9824 31136
rect 16212 31084 16264 31136
rect 16764 31127 16816 31136
rect 16764 31093 16773 31127
rect 16773 31093 16807 31127
rect 16807 31093 16816 31127
rect 16764 31084 16816 31093
rect 17408 31084 17460 31136
rect 19524 31084 19576 31136
rect 24952 31220 25004 31272
rect 26148 31084 26200 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 11244 30923 11296 30932
rect 11244 30889 11253 30923
rect 11253 30889 11287 30923
rect 11287 30889 11296 30923
rect 11244 30880 11296 30889
rect 20260 30880 20312 30932
rect 15476 30812 15528 30864
rect 22008 30880 22060 30932
rect 22836 30923 22888 30932
rect 22836 30889 22845 30923
rect 22845 30889 22879 30923
rect 22879 30889 22888 30923
rect 22836 30880 22888 30889
rect 25228 30923 25280 30932
rect 25228 30889 25237 30923
rect 25237 30889 25271 30923
rect 25271 30889 25280 30923
rect 25228 30880 25280 30889
rect 23940 30812 23992 30864
rect 25964 30812 26016 30864
rect 16488 30787 16540 30796
rect 16488 30753 16497 30787
rect 16497 30753 16531 30787
rect 16531 30753 16540 30787
rect 16488 30744 16540 30753
rect 17132 30787 17184 30796
rect 17132 30753 17141 30787
rect 17141 30753 17175 30787
rect 17175 30753 17184 30787
rect 17132 30744 17184 30753
rect 17408 30787 17460 30796
rect 17408 30753 17417 30787
rect 17417 30753 17451 30787
rect 17451 30753 17460 30787
rect 17408 30744 17460 30753
rect 10140 30676 10192 30728
rect 11796 30676 11848 30728
rect 15200 30676 15252 30728
rect 16764 30676 16816 30728
rect 20628 30744 20680 30796
rect 22836 30744 22888 30796
rect 19708 30676 19760 30728
rect 22652 30676 22704 30728
rect 12716 30608 12768 30660
rect 11060 30540 11112 30592
rect 12900 30540 12952 30592
rect 13820 30583 13872 30592
rect 13820 30549 13829 30583
rect 13829 30549 13863 30583
rect 13863 30549 13872 30583
rect 13820 30540 13872 30549
rect 14372 30608 14424 30660
rect 15844 30608 15896 30660
rect 16672 30608 16724 30660
rect 18696 30608 18748 30660
rect 21824 30608 21876 30660
rect 15384 30540 15436 30592
rect 15752 30540 15804 30592
rect 18420 30540 18472 30592
rect 20352 30540 20404 30592
rect 20812 30540 20864 30592
rect 21180 30540 21232 30592
rect 24400 30540 24452 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 11704 30336 11756 30388
rect 9680 30311 9732 30320
rect 9680 30277 9689 30311
rect 9689 30277 9723 30311
rect 9723 30277 9732 30311
rect 9680 30268 9732 30277
rect 11796 30268 11848 30320
rect 12900 30311 12952 30320
rect 12900 30277 12909 30311
rect 12909 30277 12943 30311
rect 12943 30277 12952 30311
rect 12900 30268 12952 30277
rect 13544 30336 13596 30388
rect 14556 30336 14608 30388
rect 16488 30336 16540 30388
rect 16948 30268 17000 30320
rect 21824 30336 21876 30388
rect 22284 30336 22336 30388
rect 17868 30268 17920 30320
rect 19064 30268 19116 30320
rect 20168 30268 20220 30320
rect 20996 30268 21048 30320
rect 10232 30200 10284 30252
rect 10508 30243 10560 30252
rect 10508 30209 10517 30243
rect 10517 30209 10551 30243
rect 10551 30209 10560 30243
rect 10508 30200 10560 30209
rect 15752 30200 15804 30252
rect 16304 30200 16356 30252
rect 16488 30200 16540 30252
rect 12624 30175 12676 30184
rect 12624 30141 12633 30175
rect 12633 30141 12667 30175
rect 12667 30141 12676 30175
rect 12624 30132 12676 30141
rect 14188 30132 14240 30184
rect 17040 30132 17092 30184
rect 15752 30064 15804 30116
rect 17224 30064 17276 30116
rect 18880 30200 18932 30252
rect 18972 30200 19024 30252
rect 19616 30200 19668 30252
rect 18328 30132 18380 30184
rect 19800 30132 19852 30184
rect 20444 30175 20496 30184
rect 20444 30141 20453 30175
rect 20453 30141 20487 30175
rect 20487 30141 20496 30175
rect 20444 30132 20496 30141
rect 18972 30064 19024 30116
rect 21732 30064 21784 30116
rect 15568 29996 15620 30048
rect 16764 29996 16816 30048
rect 17500 29996 17552 30048
rect 19156 29996 19208 30048
rect 19340 29996 19392 30048
rect 20168 29996 20220 30048
rect 24124 30200 24176 30252
rect 22744 30175 22796 30184
rect 22744 30141 22753 30175
rect 22753 30141 22787 30175
rect 22787 30141 22796 30175
rect 22744 30132 22796 30141
rect 23664 30132 23716 30184
rect 24952 30175 25004 30184
rect 24952 30141 24961 30175
rect 24961 30141 24995 30175
rect 24995 30141 25004 30175
rect 24952 30132 25004 30141
rect 22560 30064 22612 30116
rect 24492 30039 24544 30048
rect 24492 30005 24501 30039
rect 24501 30005 24535 30039
rect 24535 30005 24544 30039
rect 24492 29996 24544 30005
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 13820 29792 13872 29844
rect 23388 29792 23440 29844
rect 18512 29724 18564 29776
rect 19340 29724 19392 29776
rect 20352 29724 20404 29776
rect 11060 29656 11112 29708
rect 10876 29588 10928 29640
rect 12532 29656 12584 29708
rect 14188 29656 14240 29708
rect 15292 29656 15344 29708
rect 16120 29656 16172 29708
rect 16856 29656 16908 29708
rect 16948 29656 17000 29708
rect 19156 29656 19208 29708
rect 20904 29656 20956 29708
rect 13820 29588 13872 29640
rect 11520 29563 11572 29572
rect 11520 29529 11529 29563
rect 11529 29529 11563 29563
rect 11563 29529 11572 29563
rect 11520 29520 11572 29529
rect 11796 29520 11848 29572
rect 15016 29588 15068 29640
rect 16304 29588 16356 29640
rect 17132 29631 17184 29640
rect 17132 29597 17141 29631
rect 17141 29597 17175 29631
rect 17175 29597 17184 29631
rect 17132 29588 17184 29597
rect 19800 29631 19852 29640
rect 19800 29597 19809 29631
rect 19809 29597 19843 29631
rect 19843 29597 19852 29631
rect 19800 29588 19852 29597
rect 20720 29588 20772 29640
rect 21088 29699 21140 29708
rect 21088 29665 21097 29699
rect 21097 29665 21131 29699
rect 21131 29665 21140 29699
rect 21088 29656 21140 29665
rect 17316 29520 17368 29572
rect 17408 29563 17460 29572
rect 17408 29529 17417 29563
rect 17417 29529 17451 29563
rect 17451 29529 17460 29563
rect 17408 29520 17460 29529
rect 18420 29520 18472 29572
rect 19340 29520 19392 29572
rect 11888 29452 11940 29504
rect 12992 29495 13044 29504
rect 12992 29461 13001 29495
rect 13001 29461 13035 29495
rect 13035 29461 13044 29495
rect 12992 29452 13044 29461
rect 13544 29495 13596 29504
rect 13544 29461 13553 29495
rect 13553 29461 13587 29495
rect 13587 29461 13596 29495
rect 13544 29452 13596 29461
rect 14556 29452 14608 29504
rect 15292 29452 15344 29504
rect 15752 29452 15804 29504
rect 15936 29452 15988 29504
rect 16304 29452 16356 29504
rect 18328 29452 18380 29504
rect 18880 29495 18932 29504
rect 18880 29461 18889 29495
rect 18889 29461 18923 29495
rect 18923 29461 18932 29495
rect 18880 29452 18932 29461
rect 19616 29452 19668 29504
rect 20628 29495 20680 29504
rect 20628 29461 20637 29495
rect 20637 29461 20671 29495
rect 20671 29461 20680 29495
rect 20628 29452 20680 29461
rect 22836 29724 22888 29776
rect 21456 29588 21508 29640
rect 21916 29631 21968 29640
rect 21916 29597 21925 29631
rect 21925 29597 21959 29631
rect 21959 29597 21968 29631
rect 21916 29588 21968 29597
rect 24860 29656 24912 29708
rect 23756 29588 23808 29640
rect 22100 29520 22152 29572
rect 22744 29520 22796 29572
rect 23572 29452 23624 29504
rect 25228 29495 25280 29504
rect 25228 29461 25237 29495
rect 25237 29461 25271 29495
rect 25271 29461 25280 29495
rect 25228 29452 25280 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 11520 29248 11572 29300
rect 15108 29291 15160 29300
rect 15108 29257 15117 29291
rect 15117 29257 15151 29291
rect 15151 29257 15160 29291
rect 15108 29248 15160 29257
rect 15568 29248 15620 29300
rect 16856 29248 16908 29300
rect 20536 29248 20588 29300
rect 22468 29291 22520 29300
rect 22468 29257 22477 29291
rect 22477 29257 22511 29291
rect 22511 29257 22520 29291
rect 22468 29248 22520 29257
rect 24124 29248 24176 29300
rect 25780 29248 25832 29300
rect 9772 29180 9824 29232
rect 11704 29223 11756 29232
rect 11704 29189 11713 29223
rect 11713 29189 11747 29223
rect 11747 29189 11756 29223
rect 11704 29180 11756 29189
rect 13820 29180 13872 29232
rect 15936 29180 15988 29232
rect 17408 29180 17460 29232
rect 24952 29180 25004 29232
rect 11888 29112 11940 29164
rect 12624 29112 12676 29164
rect 16212 29112 16264 29164
rect 9404 29087 9456 29096
rect 9404 29053 9413 29087
rect 9413 29053 9447 29087
rect 9447 29053 9456 29087
rect 9404 29044 9456 29053
rect 14004 29044 14056 29096
rect 15660 29044 15712 29096
rect 11152 29019 11204 29028
rect 11152 28985 11161 29019
rect 11161 28985 11195 29019
rect 11195 28985 11204 29019
rect 11152 28976 11204 28985
rect 16120 29087 16172 29096
rect 16120 29053 16129 29087
rect 16129 29053 16163 29087
rect 16163 29053 16172 29087
rect 16120 29044 16172 29053
rect 16396 29044 16448 29096
rect 15476 28951 15528 28960
rect 15476 28917 15485 28951
rect 15485 28917 15519 28951
rect 15519 28917 15528 28951
rect 15476 28908 15528 28917
rect 16488 28976 16540 29028
rect 18696 29112 18748 29164
rect 20720 29112 20772 29164
rect 20812 29155 20864 29164
rect 20812 29121 20821 29155
rect 20821 29121 20855 29155
rect 20855 29121 20864 29155
rect 20812 29112 20864 29121
rect 22836 29112 22888 29164
rect 17960 28976 18012 29028
rect 17776 28908 17828 28960
rect 21180 29044 21232 29096
rect 23388 29044 23440 29096
rect 23572 29155 23624 29164
rect 23572 29121 23581 29155
rect 23581 29121 23615 29155
rect 23615 29121 23624 29155
rect 23572 29112 23624 29121
rect 24400 29155 24452 29164
rect 24400 29121 24409 29155
rect 24409 29121 24443 29155
rect 24443 29121 24452 29155
rect 24400 29112 24452 29121
rect 23940 29044 23992 29096
rect 24584 29044 24636 29096
rect 18236 28976 18288 29028
rect 18328 28976 18380 29028
rect 18696 28976 18748 29028
rect 22008 29019 22060 29028
rect 22008 28985 22017 29019
rect 22017 28985 22051 29019
rect 22051 28985 22060 29019
rect 22008 28976 22060 28985
rect 23204 29019 23256 29028
rect 23204 28985 23213 29019
rect 23213 28985 23247 29019
rect 23247 28985 23256 29019
rect 23204 28976 23256 28985
rect 23296 28976 23348 29028
rect 19248 28908 19300 28960
rect 19892 28908 19944 28960
rect 22468 28908 22520 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 8852 28704 8904 28756
rect 12716 28704 12768 28756
rect 10692 28636 10744 28688
rect 10232 28611 10284 28620
rect 10232 28577 10241 28611
rect 10241 28577 10275 28611
rect 10275 28577 10284 28611
rect 10232 28568 10284 28577
rect 11428 28568 11480 28620
rect 14924 28704 14976 28756
rect 8668 28500 8720 28552
rect 9404 28500 9456 28552
rect 11060 28543 11112 28552
rect 11060 28509 11069 28543
rect 11069 28509 11103 28543
rect 11103 28509 11112 28543
rect 11060 28500 11112 28509
rect 22376 28704 22428 28756
rect 14740 28611 14792 28620
rect 14740 28577 14749 28611
rect 14749 28577 14783 28611
rect 14783 28577 14792 28611
rect 14740 28568 14792 28577
rect 13912 28500 13964 28552
rect 14464 28500 14516 28552
rect 15936 28611 15988 28620
rect 15936 28577 15945 28611
rect 15945 28577 15979 28611
rect 15979 28577 15988 28611
rect 15936 28568 15988 28577
rect 16028 28611 16080 28620
rect 16028 28577 16037 28611
rect 16037 28577 16071 28611
rect 16071 28577 16080 28611
rect 16028 28568 16080 28577
rect 16856 28568 16908 28620
rect 17316 28568 17368 28620
rect 23020 28636 23072 28688
rect 18788 28568 18840 28620
rect 21180 28568 21232 28620
rect 23940 28704 23992 28756
rect 24124 28747 24176 28756
rect 24124 28713 24133 28747
rect 24133 28713 24167 28747
rect 24167 28713 24176 28747
rect 24124 28704 24176 28713
rect 10508 28432 10560 28484
rect 11336 28475 11388 28484
rect 11336 28441 11345 28475
rect 11345 28441 11379 28475
rect 11379 28441 11388 28475
rect 11336 28432 11388 28441
rect 9956 28364 10008 28416
rect 10416 28364 10468 28416
rect 11796 28432 11848 28484
rect 13452 28432 13504 28484
rect 15476 28432 15528 28484
rect 16672 28500 16724 28552
rect 13636 28364 13688 28416
rect 16580 28364 16632 28416
rect 16672 28407 16724 28416
rect 16672 28373 16681 28407
rect 16681 28373 16715 28407
rect 16715 28373 16724 28407
rect 16672 28364 16724 28373
rect 17776 28500 17828 28552
rect 19524 28500 19576 28552
rect 22468 28500 22520 28552
rect 23572 28500 23624 28552
rect 16948 28432 17000 28484
rect 18604 28432 18656 28484
rect 20168 28475 20220 28484
rect 20168 28441 20177 28475
rect 20177 28441 20211 28475
rect 20211 28441 20220 28475
rect 20168 28432 20220 28441
rect 20444 28432 20496 28484
rect 21916 28432 21968 28484
rect 17316 28364 17368 28416
rect 22192 28407 22244 28416
rect 22192 28373 22201 28407
rect 22201 28373 22235 28407
rect 22235 28373 22244 28407
rect 22192 28364 22244 28373
rect 24400 28432 24452 28484
rect 25780 28432 25832 28484
rect 23756 28364 23808 28416
rect 24768 28364 24820 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 10232 28160 10284 28212
rect 11704 28160 11756 28212
rect 14648 28160 14700 28212
rect 8668 28067 8720 28076
rect 8668 28033 8677 28067
rect 8677 28033 8711 28067
rect 8711 28033 8720 28067
rect 8668 28024 8720 28033
rect 11060 28024 11112 28076
rect 14372 28092 14424 28144
rect 15292 28092 15344 28144
rect 16856 28160 16908 28212
rect 16948 28203 17000 28212
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 19340 28203 19392 28212
rect 19340 28169 19349 28203
rect 19349 28169 19383 28203
rect 19383 28169 19392 28203
rect 19340 28160 19392 28169
rect 20812 28160 20864 28212
rect 25044 28160 25096 28212
rect 17868 28092 17920 28144
rect 18420 28092 18472 28144
rect 22284 28092 22336 28144
rect 8944 27999 8996 28008
rect 8944 27965 8953 27999
rect 8953 27965 8987 27999
rect 8987 27965 8996 27999
rect 8944 27956 8996 27965
rect 12440 27956 12492 28008
rect 17040 28024 17092 28076
rect 20904 28024 20956 28076
rect 21272 28024 21324 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 24216 28024 24268 28076
rect 13728 27820 13780 27872
rect 14924 27956 14976 28008
rect 15476 27820 15528 27872
rect 15752 27820 15804 27872
rect 16120 27863 16172 27872
rect 16120 27829 16129 27863
rect 16129 27829 16163 27863
rect 16163 27829 16172 27863
rect 16120 27820 16172 27829
rect 16488 27820 16540 27872
rect 20076 27956 20128 28008
rect 21088 27956 21140 28008
rect 22744 27956 22796 28008
rect 25136 27999 25188 28008
rect 25136 27965 25145 27999
rect 25145 27965 25179 27999
rect 25179 27965 25188 27999
rect 25136 27956 25188 27965
rect 19248 27888 19300 27940
rect 24584 27931 24636 27940
rect 24584 27897 24593 27931
rect 24593 27897 24627 27931
rect 24627 27897 24636 27931
rect 24584 27888 24636 27897
rect 21916 27820 21968 27872
rect 23020 27820 23072 27872
rect 23388 27820 23440 27872
rect 23572 27820 23624 27872
rect 24032 27820 24084 27872
rect 24768 27820 24820 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 10324 27616 10376 27668
rect 11704 27616 11756 27668
rect 13728 27591 13780 27600
rect 13728 27557 13737 27591
rect 13737 27557 13771 27591
rect 13771 27557 13780 27591
rect 13728 27548 13780 27557
rect 16488 27616 16540 27668
rect 18604 27659 18656 27668
rect 18604 27625 18613 27659
rect 18613 27625 18647 27659
rect 18647 27625 18656 27659
rect 18604 27616 18656 27625
rect 15292 27548 15344 27600
rect 10876 27480 10928 27532
rect 11704 27344 11756 27396
rect 15108 27412 15160 27464
rect 15292 27412 15344 27464
rect 15936 27480 15988 27532
rect 16856 27480 16908 27532
rect 14004 27344 14056 27396
rect 9312 27276 9364 27328
rect 11612 27319 11664 27328
rect 11612 27285 11621 27319
rect 11621 27285 11655 27319
rect 11655 27285 11664 27319
rect 11612 27276 11664 27285
rect 13728 27276 13780 27328
rect 14740 27276 14792 27328
rect 14832 27319 14884 27328
rect 14832 27285 14841 27319
rect 14841 27285 14875 27319
rect 14875 27285 14884 27319
rect 14832 27276 14884 27285
rect 16764 27412 16816 27464
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 19248 27480 19300 27532
rect 15752 27344 15804 27396
rect 16212 27344 16264 27396
rect 18604 27412 18656 27464
rect 16304 27276 16356 27328
rect 16488 27319 16540 27328
rect 16488 27285 16497 27319
rect 16497 27285 16531 27319
rect 16531 27285 16540 27319
rect 16488 27276 16540 27285
rect 16580 27276 16632 27328
rect 18788 27276 18840 27328
rect 23296 27616 23348 27668
rect 23480 27616 23532 27668
rect 23756 27616 23808 27668
rect 20076 27591 20128 27600
rect 20076 27557 20085 27591
rect 20085 27557 20119 27591
rect 20119 27557 20128 27591
rect 20076 27548 20128 27557
rect 21916 27548 21968 27600
rect 19708 27480 19760 27532
rect 20444 27412 20496 27464
rect 22284 27276 22336 27328
rect 22928 27344 22980 27396
rect 24492 27480 24544 27532
rect 23848 27412 23900 27464
rect 24308 27412 24360 27464
rect 22836 27319 22888 27328
rect 22836 27285 22845 27319
rect 22845 27285 22879 27319
rect 22879 27285 22888 27319
rect 22836 27276 22888 27285
rect 24124 27319 24176 27328
rect 24124 27285 24133 27319
rect 24133 27285 24167 27319
rect 24167 27285 24176 27319
rect 24124 27276 24176 27285
rect 24216 27276 24268 27328
rect 24952 27319 25004 27328
rect 24952 27285 24961 27319
rect 24961 27285 24995 27319
rect 24995 27285 25004 27319
rect 24952 27276 25004 27285
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 11336 27072 11388 27124
rect 12440 27072 12492 27124
rect 10232 27004 10284 27056
rect 13452 27047 13504 27056
rect 13452 27013 13461 27047
rect 13461 27013 13495 27047
rect 13495 27013 13504 27047
rect 13452 27004 13504 27013
rect 13912 27004 13964 27056
rect 15752 27004 15804 27056
rect 9312 26936 9364 26988
rect 9404 26979 9456 26988
rect 9404 26945 9413 26979
rect 9413 26945 9447 26979
rect 9447 26945 9456 26979
rect 9404 26936 9456 26945
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10508 26936 10560 26945
rect 12072 26936 12124 26988
rect 4252 26868 4304 26920
rect 10968 26868 11020 26920
rect 11152 26868 11204 26920
rect 13360 26800 13412 26852
rect 6828 26732 6880 26784
rect 9680 26732 9732 26784
rect 12256 26732 12308 26784
rect 14004 26732 14056 26784
rect 14280 26732 14332 26784
rect 15016 26936 15068 26988
rect 15476 26936 15528 26988
rect 15568 26936 15620 26988
rect 16212 27004 16264 27056
rect 19340 27072 19392 27124
rect 16488 27004 16540 27056
rect 17408 27004 17460 27056
rect 20168 27004 20220 27056
rect 16856 26979 16908 26988
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 17132 26936 17184 26988
rect 17868 26936 17920 26988
rect 20904 27115 20956 27124
rect 20904 27081 20913 27115
rect 20913 27081 20947 27115
rect 20947 27081 20956 27115
rect 20904 27072 20956 27081
rect 21088 27072 21140 27124
rect 21272 27072 21324 27124
rect 21824 27072 21876 27124
rect 22100 27072 22152 27124
rect 22468 27072 22520 27124
rect 14924 26868 14976 26920
rect 15936 26868 15988 26920
rect 21272 26868 21324 26920
rect 16764 26732 16816 26784
rect 19340 26800 19392 26852
rect 22376 27004 22428 27056
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22008 26936 22060 26945
rect 23664 27072 23716 27124
rect 24400 27004 24452 27056
rect 23664 26936 23716 26988
rect 25228 26936 25280 26988
rect 25964 26868 26016 26920
rect 18972 26732 19024 26784
rect 19064 26732 19116 26784
rect 20168 26732 20220 26784
rect 20812 26732 20864 26784
rect 21640 26732 21692 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 8944 26528 8996 26580
rect 9404 26528 9456 26580
rect 6828 26367 6880 26376
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 8484 26324 8536 26376
rect 10324 26460 10376 26512
rect 10600 26392 10652 26444
rect 13820 26528 13872 26580
rect 14924 26528 14976 26580
rect 15108 26528 15160 26580
rect 13452 26460 13504 26512
rect 13636 26460 13688 26512
rect 19340 26528 19392 26580
rect 25136 26528 25188 26580
rect 11612 26392 11664 26444
rect 10876 26324 10928 26376
rect 9496 26256 9548 26308
rect 13544 26324 13596 26376
rect 15016 26435 15068 26444
rect 15016 26401 15025 26435
rect 15025 26401 15059 26435
rect 15059 26401 15068 26435
rect 15016 26392 15068 26401
rect 18328 26460 18380 26512
rect 21180 26503 21232 26512
rect 21180 26469 21189 26503
rect 21189 26469 21223 26503
rect 21223 26469 21232 26503
rect 21180 26460 21232 26469
rect 25044 26460 25096 26512
rect 17868 26392 17920 26444
rect 19708 26392 19760 26444
rect 20444 26392 20496 26444
rect 21364 26392 21416 26444
rect 21916 26392 21968 26444
rect 22008 26392 22060 26444
rect 23296 26392 23348 26444
rect 24308 26392 24360 26444
rect 25320 26392 25372 26444
rect 16764 26367 16816 26376
rect 16764 26333 16773 26367
rect 16773 26333 16807 26367
rect 16807 26333 16816 26367
rect 16764 26324 16816 26333
rect 18696 26324 18748 26376
rect 18788 26324 18840 26376
rect 18972 26367 19024 26376
rect 18972 26333 18981 26367
rect 18981 26333 19015 26367
rect 19015 26333 19024 26367
rect 18972 26324 19024 26333
rect 20812 26324 20864 26376
rect 11520 26256 11572 26308
rect 12348 26188 12400 26240
rect 13544 26188 13596 26240
rect 13728 26188 13780 26240
rect 14924 26231 14976 26240
rect 14924 26197 14933 26231
rect 14933 26197 14967 26231
rect 14967 26197 14976 26231
rect 14924 26188 14976 26197
rect 15200 26256 15252 26308
rect 18420 26256 18472 26308
rect 15752 26188 15804 26240
rect 18604 26231 18656 26240
rect 18604 26197 18613 26231
rect 18613 26197 18647 26231
rect 18647 26197 18656 26231
rect 18604 26188 18656 26197
rect 23664 26324 23716 26376
rect 24400 26324 24452 26376
rect 22008 26256 22060 26308
rect 25412 26324 25464 26376
rect 25780 26256 25832 26308
rect 22100 26188 22152 26240
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 11336 25984 11388 26036
rect 12624 25984 12676 26036
rect 9680 25959 9732 25968
rect 9680 25925 9689 25959
rect 9689 25925 9723 25959
rect 9723 25925 9732 25959
rect 9680 25916 9732 25925
rect 10968 25916 11020 25968
rect 12532 25916 12584 25968
rect 13728 25984 13780 26036
rect 15384 26027 15436 26036
rect 15384 25993 15393 26027
rect 15393 25993 15427 26027
rect 15427 25993 15436 26027
rect 15384 25984 15436 25993
rect 16672 25984 16724 26036
rect 17592 25984 17644 26036
rect 18420 26027 18472 26036
rect 18420 25993 18429 26027
rect 18429 25993 18463 26027
rect 18463 25993 18472 26027
rect 18420 25984 18472 25993
rect 20628 25984 20680 26036
rect 21272 26027 21324 26036
rect 21272 25993 21281 26027
rect 21281 25993 21315 26027
rect 21315 25993 21324 26027
rect 21272 25984 21324 25993
rect 21548 26027 21600 26036
rect 21548 25993 21557 26027
rect 21557 25993 21591 26027
rect 21591 25993 21600 26027
rect 21548 25984 21600 25993
rect 22100 25984 22152 26036
rect 24124 25984 24176 26036
rect 10784 25848 10836 25900
rect 11336 25848 11388 25900
rect 11612 25848 11664 25900
rect 14924 25848 14976 25900
rect 15108 25848 15160 25900
rect 10324 25780 10376 25832
rect 10692 25780 10744 25832
rect 15476 25780 15528 25832
rect 16120 25891 16172 25900
rect 16120 25857 16129 25891
rect 16129 25857 16163 25891
rect 16163 25857 16172 25891
rect 16120 25848 16172 25857
rect 7472 25644 7524 25696
rect 8944 25687 8996 25696
rect 8944 25653 8953 25687
rect 8953 25653 8987 25687
rect 8987 25653 8996 25687
rect 8944 25644 8996 25653
rect 9036 25644 9088 25696
rect 12808 25712 12860 25764
rect 16672 25780 16724 25832
rect 11704 25644 11756 25696
rect 15752 25712 15804 25764
rect 18788 25848 18840 25900
rect 19524 25891 19576 25900
rect 19524 25857 19533 25891
rect 19533 25857 19567 25891
rect 19567 25857 19576 25891
rect 19524 25848 19576 25857
rect 21548 25848 21600 25900
rect 23296 25916 23348 25968
rect 23388 25959 23440 25968
rect 23388 25925 23397 25959
rect 23397 25925 23431 25959
rect 23431 25925 23440 25959
rect 23388 25916 23440 25925
rect 23664 25916 23716 25968
rect 18880 25780 18932 25832
rect 23388 25780 23440 25832
rect 18052 25755 18104 25764
rect 18052 25721 18061 25755
rect 18061 25721 18095 25755
rect 18095 25721 18104 25755
rect 18052 25712 18104 25721
rect 14740 25644 14792 25696
rect 15384 25644 15436 25696
rect 16488 25644 16540 25696
rect 16580 25644 16632 25696
rect 24584 25644 24636 25696
rect 25228 25687 25280 25696
rect 25228 25653 25237 25687
rect 25237 25653 25271 25687
rect 25271 25653 25280 25687
rect 25228 25644 25280 25653
rect 25412 25687 25464 25696
rect 25412 25653 25421 25687
rect 25421 25653 25455 25687
rect 25455 25653 25464 25687
rect 25412 25644 25464 25653
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 8944 25440 8996 25492
rect 10140 25440 10192 25492
rect 10600 25440 10652 25492
rect 10508 25372 10560 25424
rect 13544 25483 13596 25492
rect 13544 25449 13553 25483
rect 13553 25449 13587 25483
rect 13587 25449 13596 25483
rect 13544 25440 13596 25449
rect 10968 25304 11020 25356
rect 14464 25304 14516 25356
rect 13452 25236 13504 25288
rect 14648 25372 14700 25424
rect 14832 25304 14884 25356
rect 15568 25304 15620 25356
rect 18696 25483 18748 25492
rect 18696 25449 18705 25483
rect 18705 25449 18739 25483
rect 18739 25449 18748 25483
rect 18696 25440 18748 25449
rect 19156 25440 19208 25492
rect 19524 25440 19576 25492
rect 20720 25440 20772 25492
rect 21916 25440 21968 25492
rect 25688 25440 25740 25492
rect 24124 25372 24176 25424
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 17592 25236 17644 25288
rect 19064 25236 19116 25288
rect 9680 25168 9732 25220
rect 10784 25168 10836 25220
rect 12624 25168 12676 25220
rect 10140 25100 10192 25152
rect 13820 25168 13872 25220
rect 14188 25168 14240 25220
rect 15016 25168 15068 25220
rect 16764 25168 16816 25220
rect 18512 25168 18564 25220
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 20996 25304 21048 25356
rect 21456 25236 21508 25288
rect 21916 25279 21968 25288
rect 21916 25245 21925 25279
rect 21925 25245 21959 25279
rect 21959 25245 21968 25279
rect 21916 25236 21968 25245
rect 22560 25236 22612 25288
rect 24400 25236 24452 25288
rect 21180 25168 21232 25220
rect 22836 25168 22888 25220
rect 24952 25168 25004 25220
rect 13176 25100 13228 25152
rect 13912 25100 13964 25152
rect 14648 25100 14700 25152
rect 16028 25143 16080 25152
rect 16028 25109 16037 25143
rect 16037 25109 16071 25143
rect 16071 25109 16080 25143
rect 16028 25100 16080 25109
rect 16396 25100 16448 25152
rect 18328 25100 18380 25152
rect 20812 25143 20864 25152
rect 20812 25109 20821 25143
rect 20821 25109 20855 25143
rect 20855 25109 20864 25143
rect 20812 25100 20864 25109
rect 20904 25100 20956 25152
rect 21916 25100 21968 25152
rect 22560 25100 22612 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 9588 24896 9640 24948
rect 10508 24896 10560 24948
rect 15384 24896 15436 24948
rect 16120 24896 16172 24948
rect 16304 24896 16356 24948
rect 16488 24896 16540 24948
rect 17500 24896 17552 24948
rect 10784 24828 10836 24880
rect 12808 24828 12860 24880
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 8576 24803 8628 24812
rect 8576 24769 8585 24803
rect 8585 24769 8619 24803
rect 8619 24769 8628 24803
rect 8576 24760 8628 24769
rect 11704 24803 11756 24812
rect 11704 24769 11713 24803
rect 11713 24769 11747 24803
rect 11747 24769 11756 24803
rect 11704 24760 11756 24769
rect 13176 24803 13228 24812
rect 13176 24769 13185 24803
rect 13185 24769 13219 24803
rect 13219 24769 13228 24803
rect 13176 24760 13228 24769
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13544 24828 13596 24880
rect 13728 24828 13780 24880
rect 15660 24828 15712 24880
rect 17684 24896 17736 24948
rect 18604 24896 18656 24948
rect 19156 24896 19208 24948
rect 20720 24896 20772 24948
rect 24032 24896 24084 24948
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 15476 24760 15528 24812
rect 16212 24760 16264 24812
rect 18696 24828 18748 24880
rect 19984 24828 20036 24880
rect 21916 24828 21968 24880
rect 25228 24828 25280 24880
rect 15016 24692 15068 24744
rect 16488 24692 16540 24744
rect 17316 24692 17368 24744
rect 19340 24760 19392 24812
rect 19708 24803 19760 24812
rect 19708 24769 19717 24803
rect 19717 24769 19751 24803
rect 19751 24769 19760 24803
rect 19708 24760 19760 24769
rect 21272 24760 21324 24812
rect 18328 24692 18380 24744
rect 9864 24556 9916 24608
rect 10692 24556 10744 24608
rect 10876 24556 10928 24608
rect 12532 24556 12584 24608
rect 13360 24556 13412 24608
rect 18420 24624 18472 24676
rect 18512 24667 18564 24676
rect 18512 24633 18521 24667
rect 18521 24633 18555 24667
rect 18555 24633 18564 24667
rect 18512 24624 18564 24633
rect 16488 24556 16540 24608
rect 16948 24556 17000 24608
rect 19064 24735 19116 24744
rect 19064 24701 19073 24735
rect 19073 24701 19107 24735
rect 19107 24701 19116 24735
rect 19064 24692 19116 24701
rect 21364 24692 21416 24744
rect 22192 24624 22244 24676
rect 22652 24692 22704 24744
rect 23296 24692 23348 24744
rect 23940 24692 23992 24744
rect 21272 24556 21324 24608
rect 22100 24599 22152 24608
rect 22100 24565 22109 24599
rect 22109 24565 22143 24599
rect 22143 24565 22152 24599
rect 22100 24556 22152 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 25228 24556 25280 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 10048 24395 10100 24404
rect 10048 24361 10057 24395
rect 10057 24361 10091 24395
rect 10091 24361 10100 24395
rect 10048 24352 10100 24361
rect 6460 24148 6512 24200
rect 9588 24148 9640 24200
rect 14648 24352 14700 24404
rect 15660 24352 15712 24404
rect 14464 24284 14516 24336
rect 10876 24216 10928 24268
rect 11520 24259 11572 24268
rect 11520 24225 11529 24259
rect 11529 24225 11563 24259
rect 11563 24225 11572 24259
rect 11520 24216 11572 24225
rect 20260 24352 20312 24404
rect 21548 24395 21600 24404
rect 21548 24361 21557 24395
rect 21557 24361 21591 24395
rect 21591 24361 21600 24395
rect 21548 24352 21600 24361
rect 25136 24352 25188 24404
rect 17132 24284 17184 24336
rect 19708 24284 19760 24336
rect 11244 24191 11296 24200
rect 11244 24157 11253 24191
rect 11253 24157 11287 24191
rect 11287 24157 11296 24191
rect 11244 24148 11296 24157
rect 12624 24148 12676 24200
rect 13084 24148 13136 24200
rect 17040 24216 17092 24268
rect 18880 24216 18932 24268
rect 15384 24148 15436 24200
rect 17500 24148 17552 24200
rect 18420 24148 18472 24200
rect 20996 24216 21048 24268
rect 6920 24012 6972 24064
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 10508 24055 10560 24064
rect 10508 24021 10517 24055
rect 10517 24021 10551 24055
rect 10551 24021 10560 24055
rect 10508 24012 10560 24021
rect 20444 24123 20496 24132
rect 20444 24089 20453 24123
rect 20453 24089 20487 24123
rect 20487 24089 20496 24123
rect 20444 24080 20496 24089
rect 20720 24148 20772 24200
rect 21640 24148 21692 24200
rect 21916 24148 21968 24200
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 21272 24080 21324 24132
rect 22284 24123 22336 24132
rect 22284 24089 22293 24123
rect 22293 24089 22327 24123
rect 22327 24089 22336 24123
rect 22284 24080 22336 24089
rect 23664 24080 23716 24132
rect 25320 24080 25372 24132
rect 13452 24012 13504 24064
rect 13728 24012 13780 24064
rect 13912 24012 13964 24064
rect 16672 24012 16724 24064
rect 17224 24055 17276 24064
rect 17224 24021 17233 24055
rect 17233 24021 17267 24055
rect 17267 24021 17276 24055
rect 17224 24012 17276 24021
rect 18420 24012 18472 24064
rect 18512 24055 18564 24064
rect 18512 24021 18521 24055
rect 18521 24021 18555 24055
rect 18555 24021 18564 24055
rect 18512 24012 18564 24021
rect 18788 24012 18840 24064
rect 19156 24012 19208 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 19892 24055 19944 24064
rect 19892 24021 19901 24055
rect 19901 24021 19935 24055
rect 19935 24021 19944 24055
rect 19892 24012 19944 24021
rect 20352 24012 20404 24064
rect 23848 24012 23900 24064
rect 24032 24055 24084 24064
rect 24032 24021 24041 24055
rect 24041 24021 24075 24055
rect 24075 24021 24084 24055
rect 24032 24012 24084 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 6460 23851 6512 23860
rect 6460 23817 6469 23851
rect 6469 23817 6503 23851
rect 6503 23817 6512 23851
rect 6460 23808 6512 23817
rect 9128 23851 9180 23860
rect 9128 23817 9137 23851
rect 9137 23817 9171 23851
rect 9171 23817 9180 23851
rect 9128 23808 9180 23817
rect 10048 23808 10100 23860
rect 10324 23808 10376 23860
rect 7656 23740 7708 23792
rect 13084 23851 13136 23860
rect 13084 23817 13093 23851
rect 13093 23817 13127 23851
rect 13127 23817 13136 23851
rect 13084 23808 13136 23817
rect 13912 23851 13964 23860
rect 13912 23817 13921 23851
rect 13921 23817 13955 23851
rect 13955 23817 13964 23851
rect 13912 23808 13964 23817
rect 16028 23808 16080 23860
rect 18512 23808 18564 23860
rect 19248 23808 19300 23860
rect 12072 23740 12124 23792
rect 6920 23715 6972 23724
rect 6920 23681 6929 23715
rect 6929 23681 6963 23715
rect 6963 23681 6972 23715
rect 6920 23672 6972 23681
rect 10324 23672 10376 23724
rect 14004 23783 14056 23792
rect 14004 23749 14013 23783
rect 14013 23749 14047 23783
rect 14047 23749 14056 23783
rect 14004 23740 14056 23749
rect 19524 23808 19576 23860
rect 19708 23808 19760 23860
rect 24216 23808 24268 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 25412 23808 25464 23860
rect 7196 23647 7248 23656
rect 7196 23613 7205 23647
rect 7205 23613 7239 23647
rect 7239 23613 7248 23647
rect 7196 23604 7248 23613
rect 9680 23647 9732 23656
rect 9680 23613 9689 23647
rect 9689 23613 9723 23647
rect 9723 23613 9732 23647
rect 9680 23604 9732 23613
rect 10140 23604 10192 23656
rect 12808 23604 12860 23656
rect 13268 23536 13320 23588
rect 8392 23468 8444 23520
rect 12624 23468 12676 23520
rect 14648 23672 14700 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 19064 23715 19116 23724
rect 19064 23681 19073 23715
rect 19073 23681 19107 23715
rect 19107 23681 19116 23715
rect 19064 23672 19116 23681
rect 20076 23604 20128 23656
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 21456 23672 21508 23681
rect 21824 23672 21876 23724
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 23388 23740 23440 23792
rect 25320 23783 25372 23792
rect 25320 23749 25329 23783
rect 25329 23749 25363 23783
rect 25363 23749 25372 23783
rect 25320 23740 25372 23749
rect 22652 23604 22704 23613
rect 23204 23647 23256 23656
rect 23204 23613 23213 23647
rect 23213 23613 23247 23647
rect 23247 23613 23256 23647
rect 23204 23604 23256 23613
rect 25688 23604 25740 23656
rect 21456 23536 21508 23588
rect 21916 23536 21968 23588
rect 15476 23468 15528 23520
rect 20628 23468 20680 23520
rect 21088 23468 21140 23520
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 22008 23511 22060 23520
rect 22008 23477 22017 23511
rect 22017 23477 22051 23511
rect 22051 23477 22060 23511
rect 22008 23468 22060 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 8484 23264 8536 23316
rect 12808 23264 12860 23316
rect 21548 23264 21600 23316
rect 21824 23264 21876 23316
rect 23664 23264 23716 23316
rect 7656 23128 7708 23180
rect 6276 23103 6328 23112
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 16488 23196 16540 23248
rect 7840 23128 7892 23180
rect 9404 23128 9456 23180
rect 10692 23128 10744 23180
rect 13452 23128 13504 23180
rect 15200 23128 15252 23180
rect 15936 23128 15988 23180
rect 12532 23060 12584 23112
rect 9680 22992 9732 23044
rect 10784 22992 10836 23044
rect 10876 22967 10928 22976
rect 10876 22933 10885 22967
rect 10885 22933 10919 22967
rect 10919 22933 10928 22967
rect 10876 22924 10928 22933
rect 12164 22924 12216 22976
rect 14280 23103 14332 23112
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 21640 23196 21692 23248
rect 18604 23128 18656 23180
rect 19340 23171 19392 23180
rect 19340 23137 19349 23171
rect 19349 23137 19383 23171
rect 19383 23137 19392 23171
rect 19340 23128 19392 23137
rect 19616 23128 19668 23180
rect 19892 23128 19944 23180
rect 20720 23128 20772 23180
rect 20812 23128 20864 23180
rect 24492 23128 24544 23180
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 20168 23060 20220 23112
rect 20260 23103 20312 23112
rect 20260 23069 20269 23103
rect 20269 23069 20303 23103
rect 20303 23069 20312 23103
rect 20260 23060 20312 23069
rect 20628 23060 20680 23112
rect 21824 23060 21876 23112
rect 25596 23060 25648 23112
rect 14740 22924 14792 22976
rect 15016 22992 15068 23044
rect 23388 22992 23440 23044
rect 25780 22992 25832 23044
rect 26148 22992 26200 23044
rect 15844 22924 15896 22976
rect 16120 22924 16172 22976
rect 16488 22967 16540 22976
rect 16488 22933 16497 22967
rect 16497 22933 16531 22967
rect 16531 22933 16540 22967
rect 16488 22924 16540 22933
rect 16672 22924 16724 22976
rect 17868 22924 17920 22976
rect 18788 22924 18840 22976
rect 19616 22924 19668 22976
rect 19892 22967 19944 22976
rect 19892 22933 19901 22967
rect 19901 22933 19935 22967
rect 19935 22933 19944 22967
rect 19892 22924 19944 22933
rect 20720 22924 20772 22976
rect 24676 22924 24728 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 12348 22720 12400 22772
rect 9128 22652 9180 22704
rect 10140 22652 10192 22704
rect 10784 22652 10836 22704
rect 13360 22652 13412 22704
rect 7196 22584 7248 22636
rect 7840 22584 7892 22636
rect 14924 22720 14976 22772
rect 16212 22720 16264 22772
rect 16856 22720 16908 22772
rect 18696 22720 18748 22772
rect 19156 22763 19208 22772
rect 19156 22729 19165 22763
rect 19165 22729 19199 22763
rect 19199 22729 19208 22763
rect 19156 22720 19208 22729
rect 19432 22720 19484 22772
rect 20904 22720 20956 22772
rect 21364 22763 21416 22772
rect 21364 22729 21373 22763
rect 21373 22729 21407 22763
rect 21407 22729 21416 22763
rect 21364 22720 21416 22729
rect 14740 22652 14792 22704
rect 15844 22652 15896 22704
rect 18236 22652 18288 22704
rect 18328 22695 18380 22704
rect 18328 22661 18337 22695
rect 18337 22661 18371 22695
rect 18371 22661 18380 22695
rect 18328 22652 18380 22661
rect 19064 22652 19116 22704
rect 21732 22652 21784 22704
rect 16672 22584 16724 22636
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 7656 22516 7708 22568
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 8484 22448 8536 22500
rect 7840 22380 7892 22432
rect 10692 22423 10744 22432
rect 10692 22389 10701 22423
rect 10701 22389 10735 22423
rect 10735 22389 10744 22423
rect 10692 22380 10744 22389
rect 11060 22380 11112 22432
rect 13544 22423 13596 22432
rect 13544 22389 13553 22423
rect 13553 22389 13587 22423
rect 13587 22389 13596 22423
rect 13544 22380 13596 22389
rect 15476 22516 15528 22568
rect 16396 22559 16448 22568
rect 16396 22525 16405 22559
rect 16405 22525 16439 22559
rect 16439 22525 16448 22559
rect 16396 22516 16448 22525
rect 17500 22516 17552 22568
rect 20076 22559 20128 22568
rect 20076 22525 20085 22559
rect 20085 22525 20119 22559
rect 20119 22525 20128 22559
rect 20076 22516 20128 22525
rect 24952 22584 25004 22636
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 14280 22380 14332 22432
rect 16856 22448 16908 22500
rect 20168 22448 20220 22500
rect 26056 22448 26108 22500
rect 18696 22380 18748 22432
rect 19524 22423 19576 22432
rect 19524 22389 19533 22423
rect 19533 22389 19567 22423
rect 19567 22389 19576 22423
rect 19524 22380 19576 22389
rect 25320 22380 25372 22432
rect 25596 22380 25648 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 6276 22176 6328 22228
rect 15108 22176 15160 22228
rect 19248 22219 19300 22228
rect 19248 22185 19257 22219
rect 19257 22185 19291 22219
rect 19291 22185 19300 22219
rect 19248 22176 19300 22185
rect 20168 22176 20220 22228
rect 21088 22176 21140 22228
rect 25320 22176 25372 22228
rect 10600 22108 10652 22160
rect 13360 22108 13412 22160
rect 7104 22040 7156 22092
rect 3700 21836 3752 21888
rect 8208 21972 8260 22024
rect 9588 21972 9640 22024
rect 9956 21972 10008 22024
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 13452 22040 13504 22092
rect 13820 22040 13872 22092
rect 13544 21972 13596 22024
rect 13728 21972 13780 22024
rect 16120 22040 16172 22092
rect 16580 21972 16632 22024
rect 17500 21972 17552 22024
rect 18788 21972 18840 22024
rect 19340 22040 19392 22092
rect 6736 21904 6788 21956
rect 8668 21836 8720 21888
rect 10232 21879 10284 21888
rect 10232 21845 10241 21879
rect 10241 21845 10275 21879
rect 10275 21845 10284 21879
rect 10232 21836 10284 21845
rect 10600 21879 10652 21888
rect 10600 21845 10609 21879
rect 10609 21845 10643 21879
rect 10643 21845 10652 21879
rect 10600 21836 10652 21845
rect 10784 21836 10836 21888
rect 12624 21879 12676 21888
rect 12624 21845 12633 21879
rect 12633 21845 12667 21879
rect 12667 21845 12676 21879
rect 12624 21836 12676 21845
rect 13176 21836 13228 21888
rect 14556 21836 14608 21888
rect 15108 21836 15160 21888
rect 17868 21904 17920 21956
rect 19248 21904 19300 21956
rect 20812 21972 20864 22024
rect 17776 21879 17828 21888
rect 17776 21845 17785 21879
rect 17785 21845 17819 21879
rect 17819 21845 17828 21879
rect 17776 21836 17828 21845
rect 18880 21879 18932 21888
rect 18880 21845 18889 21879
rect 18889 21845 18923 21879
rect 18923 21845 18932 21879
rect 18880 21836 18932 21845
rect 20812 21836 20864 21888
rect 21456 22083 21508 22092
rect 21456 22049 21465 22083
rect 21465 22049 21499 22083
rect 21499 22049 21508 22083
rect 21456 22040 21508 22049
rect 21732 22040 21784 22092
rect 21088 21972 21140 22024
rect 24032 22040 24084 22092
rect 24492 22040 24544 22092
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 25228 22083 25280 22092
rect 25228 22049 25237 22083
rect 25237 22049 25271 22083
rect 25271 22049 25280 22083
rect 25228 22040 25280 22049
rect 22008 21904 22060 21956
rect 21088 21879 21140 21888
rect 21088 21845 21097 21879
rect 21097 21845 21131 21879
rect 21131 21845 21140 21879
rect 21088 21836 21140 21845
rect 21180 21836 21232 21888
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 24952 21879 25004 21888
rect 24952 21845 24961 21879
rect 24961 21845 24995 21879
rect 24995 21845 25004 21879
rect 24952 21836 25004 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 8852 21632 8904 21684
rect 9680 21632 9732 21684
rect 10416 21675 10468 21684
rect 10416 21641 10425 21675
rect 10425 21641 10459 21675
rect 10459 21641 10468 21675
rect 10416 21632 10468 21641
rect 4712 21496 4764 21548
rect 8668 21564 8720 21616
rect 7472 21496 7524 21548
rect 11980 21564 12032 21616
rect 15108 21632 15160 21684
rect 12808 21564 12860 21616
rect 13176 21607 13228 21616
rect 13176 21573 13185 21607
rect 13185 21573 13219 21607
rect 13219 21573 13228 21607
rect 13176 21564 13228 21573
rect 14464 21564 14516 21616
rect 14648 21564 14700 21616
rect 16672 21632 16724 21684
rect 18604 21632 18656 21684
rect 19616 21632 19668 21684
rect 20812 21632 20864 21684
rect 21364 21632 21416 21684
rect 17132 21564 17184 21616
rect 19708 21564 19760 21616
rect 21088 21564 21140 21616
rect 21456 21564 21508 21616
rect 22192 21564 22244 21616
rect 22468 21607 22520 21616
rect 22468 21573 22477 21607
rect 22477 21573 22511 21607
rect 22511 21573 22520 21607
rect 22468 21564 22520 21573
rect 25596 21564 25648 21616
rect 10692 21360 10744 21412
rect 6828 21292 6880 21344
rect 11060 21496 11112 21548
rect 16120 21496 16172 21548
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 18972 21496 19024 21548
rect 20168 21496 20220 21548
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 20444 21496 20496 21548
rect 22008 21496 22060 21548
rect 22100 21496 22152 21548
rect 22284 21496 22336 21548
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 10876 21360 10928 21412
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 18604 21428 18656 21480
rect 19064 21428 19116 21480
rect 20812 21428 20864 21480
rect 22468 21428 22520 21480
rect 11244 21360 11296 21412
rect 12348 21360 12400 21412
rect 11612 21292 11664 21344
rect 14188 21292 14240 21344
rect 14648 21335 14700 21344
rect 14648 21301 14657 21335
rect 14657 21301 14691 21335
rect 14691 21301 14700 21335
rect 14648 21292 14700 21301
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 16396 21292 16448 21344
rect 18788 21292 18840 21344
rect 19432 21292 19484 21344
rect 20904 21292 20956 21344
rect 22284 21360 22336 21412
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 24216 21428 24268 21480
rect 24032 21292 24084 21344
rect 24492 21292 24544 21344
rect 25504 21292 25556 21344
rect 25872 21292 25924 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 10324 21088 10376 21140
rect 10692 21088 10744 21140
rect 25136 21088 25188 21140
rect 25504 21088 25556 21140
rect 7656 20884 7708 20936
rect 7840 20884 7892 20936
rect 11520 21020 11572 21072
rect 13360 21020 13412 21072
rect 13544 21020 13596 21072
rect 14924 21020 14976 21072
rect 15292 21063 15344 21072
rect 15292 21029 15301 21063
rect 15301 21029 15335 21063
rect 15335 21029 15344 21063
rect 15292 21020 15344 21029
rect 16396 21063 16448 21072
rect 16396 21029 16405 21063
rect 16405 21029 16439 21063
rect 16439 21029 16448 21063
rect 16396 21020 16448 21029
rect 18604 21063 18656 21072
rect 18604 21029 18613 21063
rect 18613 21029 18647 21063
rect 18647 21029 18656 21063
rect 18604 21020 18656 21029
rect 18972 21063 19024 21072
rect 18972 21029 18981 21063
rect 18981 21029 19015 21063
rect 19015 21029 19024 21063
rect 18972 21020 19024 21029
rect 19708 21020 19760 21072
rect 9680 20952 9732 21004
rect 11244 20952 11296 21004
rect 12624 20952 12676 21004
rect 11060 20884 11112 20936
rect 14464 20884 14516 20936
rect 16304 20952 16356 21004
rect 20352 20952 20404 21004
rect 21824 21063 21876 21072
rect 21824 21029 21833 21063
rect 21833 21029 21867 21063
rect 21867 21029 21876 21063
rect 21824 21020 21876 21029
rect 22008 21020 22060 21072
rect 24952 21020 25004 21072
rect 16764 20884 16816 20936
rect 9128 20816 9180 20868
rect 5080 20791 5132 20800
rect 5080 20757 5089 20791
rect 5089 20757 5123 20791
rect 5123 20757 5132 20791
rect 5080 20748 5132 20757
rect 6644 20748 6696 20800
rect 7472 20791 7524 20800
rect 7472 20757 7481 20791
rect 7481 20757 7515 20791
rect 7515 20757 7524 20791
rect 7472 20748 7524 20757
rect 10692 20748 10744 20800
rect 11888 20859 11940 20868
rect 11888 20825 11897 20859
rect 11897 20825 11931 20859
rect 11931 20825 11940 20859
rect 11888 20816 11940 20825
rect 14556 20816 14608 20868
rect 16304 20816 16356 20868
rect 17040 20884 17092 20936
rect 19616 20884 19668 20936
rect 25044 20952 25096 21004
rect 13360 20791 13412 20800
rect 13360 20757 13369 20791
rect 13369 20757 13403 20791
rect 13403 20757 13412 20791
rect 13360 20748 13412 20757
rect 13636 20791 13688 20800
rect 13636 20757 13645 20791
rect 13645 20757 13679 20791
rect 13679 20757 13688 20791
rect 13636 20748 13688 20757
rect 14188 20791 14240 20800
rect 14188 20757 14197 20791
rect 14197 20757 14231 20791
rect 14231 20757 14240 20791
rect 14188 20748 14240 20757
rect 19064 20816 19116 20868
rect 19156 20816 19208 20868
rect 21824 20884 21876 20936
rect 23756 20884 23808 20936
rect 23940 20884 23992 20936
rect 23112 20816 23164 20868
rect 23664 20816 23716 20868
rect 17316 20748 17368 20800
rect 17684 20748 17736 20800
rect 18604 20748 18656 20800
rect 18880 20748 18932 20800
rect 19248 20748 19300 20800
rect 20444 20748 20496 20800
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 20812 20748 20864 20800
rect 21456 20748 21508 20800
rect 21824 20748 21876 20800
rect 24584 20748 24636 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 6736 20544 6788 20596
rect 10600 20544 10652 20596
rect 11888 20544 11940 20596
rect 14648 20544 14700 20596
rect 17592 20544 17644 20596
rect 8116 20476 8168 20528
rect 10140 20476 10192 20528
rect 6000 20408 6052 20460
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 7288 20408 7340 20460
rect 11060 20408 11112 20460
rect 17500 20476 17552 20528
rect 19156 20587 19208 20596
rect 19156 20553 19165 20587
rect 19165 20553 19199 20587
rect 19199 20553 19208 20587
rect 19156 20544 19208 20553
rect 19340 20587 19392 20596
rect 19340 20553 19349 20587
rect 19349 20553 19383 20587
rect 19383 20553 19392 20587
rect 19340 20544 19392 20553
rect 21548 20544 21600 20596
rect 22376 20544 22428 20596
rect 23204 20587 23256 20596
rect 23204 20553 23213 20587
rect 23213 20553 23247 20587
rect 23247 20553 23256 20587
rect 23204 20544 23256 20553
rect 25504 20544 25556 20596
rect 5080 20340 5132 20392
rect 9128 20340 9180 20392
rect 12256 20340 12308 20392
rect 9588 20272 9640 20324
rect 16856 20408 16908 20460
rect 20720 20408 20772 20460
rect 22652 20476 22704 20528
rect 21548 20408 21600 20460
rect 13728 20340 13780 20392
rect 16396 20340 16448 20392
rect 19248 20340 19300 20392
rect 19340 20340 19392 20392
rect 20444 20340 20496 20392
rect 22284 20340 22336 20392
rect 23848 20476 23900 20528
rect 25136 20476 25188 20528
rect 23296 20408 23348 20460
rect 22008 20315 22060 20324
rect 22008 20281 22017 20315
rect 22017 20281 22051 20315
rect 22051 20281 22060 20315
rect 22008 20272 22060 20281
rect 6920 20204 6972 20256
rect 8576 20204 8628 20256
rect 12624 20204 12676 20256
rect 15016 20204 15068 20256
rect 15844 20204 15896 20256
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 17684 20204 17736 20256
rect 19616 20247 19668 20256
rect 19616 20213 19625 20247
rect 19625 20213 19659 20247
rect 19659 20213 19668 20247
rect 19616 20204 19668 20213
rect 20628 20204 20680 20256
rect 21088 20204 21140 20256
rect 21548 20204 21600 20256
rect 23848 20383 23900 20392
rect 23848 20349 23857 20383
rect 23857 20349 23891 20383
rect 23891 20349 23900 20383
rect 23848 20340 23900 20349
rect 23112 20247 23164 20256
rect 23112 20213 23121 20247
rect 23121 20213 23155 20247
rect 23155 20213 23164 20247
rect 23112 20204 23164 20213
rect 23664 20204 23716 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 7748 20000 7800 20052
rect 7932 20000 7984 20052
rect 9680 20000 9732 20052
rect 12532 20000 12584 20052
rect 12900 20000 12952 20052
rect 12440 19932 12492 19984
rect 12992 19932 13044 19984
rect 16672 20000 16724 20052
rect 16764 20000 16816 20052
rect 17500 20000 17552 20052
rect 18236 20000 18288 20052
rect 18328 20000 18380 20052
rect 18880 20000 18932 20052
rect 19800 20000 19852 20052
rect 22836 20000 22888 20052
rect 4344 19907 4396 19916
rect 4344 19873 4353 19907
rect 4353 19873 4387 19907
rect 4387 19873 4396 19907
rect 4344 19864 4396 19873
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 7748 19864 7800 19916
rect 8484 19864 8536 19916
rect 9036 19864 9088 19916
rect 6920 19796 6972 19848
rect 7288 19796 7340 19848
rect 11152 19864 11204 19916
rect 18972 19932 19024 19984
rect 19156 19932 19208 19984
rect 20628 19932 20680 19984
rect 12256 19796 12308 19848
rect 12532 19796 12584 19848
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 7196 19660 7248 19712
rect 8944 19728 8996 19780
rect 9220 19728 9272 19780
rect 14004 19796 14056 19848
rect 14464 19907 14516 19916
rect 14464 19873 14473 19907
rect 14473 19873 14507 19907
rect 14507 19873 14516 19907
rect 14464 19864 14516 19873
rect 14648 19864 14700 19916
rect 18788 19864 18840 19916
rect 15292 19796 15344 19848
rect 17500 19796 17552 19848
rect 18512 19796 18564 19848
rect 20076 19864 20128 19916
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 8852 19660 8904 19712
rect 9312 19660 9364 19712
rect 11336 19660 11388 19712
rect 11888 19660 11940 19712
rect 13636 19728 13688 19780
rect 15108 19728 15160 19780
rect 16948 19728 17000 19780
rect 19156 19728 19208 19780
rect 19340 19728 19392 19780
rect 21732 19728 21784 19780
rect 12256 19660 12308 19712
rect 13912 19660 13964 19712
rect 15568 19703 15620 19712
rect 15568 19669 15577 19703
rect 15577 19669 15611 19703
rect 15611 19669 15620 19703
rect 15568 19660 15620 19669
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 18512 19660 18564 19712
rect 19064 19660 19116 19712
rect 20352 19703 20404 19712
rect 20352 19669 20361 19703
rect 20361 19669 20395 19703
rect 20395 19669 20404 19703
rect 20352 19660 20404 19669
rect 24952 19864 25004 19916
rect 22192 19796 22244 19848
rect 24308 19796 24360 19848
rect 23388 19728 23440 19780
rect 22376 19660 22428 19712
rect 25136 19660 25188 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 4344 19456 4396 19508
rect 6000 19499 6052 19508
rect 6000 19465 6009 19499
rect 6009 19465 6043 19499
rect 6043 19465 6052 19499
rect 6000 19456 6052 19465
rect 8484 19456 8536 19508
rect 8576 19456 8628 19508
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 7840 19388 7892 19440
rect 8300 19388 8352 19440
rect 9496 19456 9548 19508
rect 9772 19388 9824 19440
rect 10416 19456 10468 19508
rect 15200 19456 15252 19508
rect 12072 19388 12124 19440
rect 7288 19363 7340 19372
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4252 19252 4304 19304
rect 6000 19184 6052 19236
rect 7932 19252 7984 19304
rect 11428 19320 11480 19372
rect 11888 19320 11940 19372
rect 12992 19388 13044 19440
rect 13544 19388 13596 19440
rect 12900 19320 12952 19372
rect 13728 19320 13780 19372
rect 17500 19499 17552 19508
rect 17500 19465 17509 19499
rect 17509 19465 17543 19499
rect 17543 19465 17552 19499
rect 17500 19456 17552 19465
rect 19340 19456 19392 19508
rect 16212 19388 16264 19440
rect 16396 19320 16448 19372
rect 18420 19320 18472 19372
rect 19064 19320 19116 19372
rect 19340 19320 19392 19372
rect 20628 19456 20680 19508
rect 20076 19388 20128 19440
rect 22284 19456 22336 19508
rect 23296 19456 23348 19508
rect 23756 19456 23808 19508
rect 24676 19499 24728 19508
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 25504 19499 25556 19508
rect 25504 19465 25513 19499
rect 25513 19465 25547 19499
rect 25547 19465 25556 19499
rect 25504 19456 25556 19465
rect 22376 19388 22428 19440
rect 8576 19184 8628 19236
rect 9312 19184 9364 19236
rect 2780 19116 2832 19168
rect 8208 19116 8260 19168
rect 10600 19159 10652 19168
rect 10600 19125 10609 19159
rect 10609 19125 10643 19159
rect 10643 19125 10652 19159
rect 10600 19116 10652 19125
rect 10876 19116 10928 19168
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 11980 19159 12032 19168
rect 11980 19125 11989 19159
rect 11989 19125 12023 19159
rect 12023 19125 12032 19159
rect 11980 19116 12032 19125
rect 13452 19295 13504 19304
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 12348 19184 12400 19236
rect 12716 19184 12768 19236
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 15108 19252 15160 19304
rect 18328 19252 18380 19304
rect 18972 19252 19024 19304
rect 22744 19252 22796 19304
rect 23940 19320 23992 19372
rect 15752 19184 15804 19236
rect 18144 19184 18196 19236
rect 18236 19184 18288 19236
rect 14188 19116 14240 19168
rect 15384 19116 15436 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 16304 19116 16356 19168
rect 19064 19116 19116 19168
rect 23480 19184 23532 19236
rect 24492 19252 24544 19304
rect 25136 19252 25188 19304
rect 26148 19252 26200 19304
rect 20076 19116 20128 19168
rect 20536 19116 20588 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 4252 18751 4304 18760
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 13912 18912 13964 18964
rect 15016 18912 15068 18964
rect 6000 18887 6052 18896
rect 6000 18853 6009 18887
rect 6009 18853 6043 18887
rect 6043 18853 6052 18887
rect 6000 18844 6052 18853
rect 9588 18887 9640 18896
rect 9588 18853 9597 18887
rect 9597 18853 9631 18887
rect 9631 18853 9640 18887
rect 9588 18844 9640 18853
rect 11336 18844 11388 18896
rect 16396 18844 16448 18896
rect 7288 18776 7340 18828
rect 6000 18708 6052 18760
rect 8116 18776 8168 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 10600 18776 10652 18828
rect 11704 18776 11756 18828
rect 12348 18776 12400 18828
rect 14464 18776 14516 18828
rect 8576 18708 8628 18760
rect 8668 18708 8720 18760
rect 11060 18708 11112 18760
rect 4068 18615 4120 18624
rect 4068 18581 4077 18615
rect 4077 18581 4111 18615
rect 4111 18581 4120 18615
rect 4068 18572 4120 18581
rect 4528 18572 4580 18624
rect 6644 18640 6696 18692
rect 12164 18640 12216 18692
rect 12256 18683 12308 18692
rect 12256 18649 12265 18683
rect 12265 18649 12299 18683
rect 12299 18649 12308 18683
rect 12256 18640 12308 18649
rect 13544 18640 13596 18692
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 11060 18572 11112 18624
rect 11336 18572 11388 18624
rect 12072 18572 12124 18624
rect 12348 18572 12400 18624
rect 13636 18572 13688 18624
rect 15200 18708 15252 18760
rect 16488 18819 16540 18828
rect 16488 18785 16497 18819
rect 16497 18785 16531 18819
rect 16531 18785 16540 18819
rect 16488 18776 16540 18785
rect 18144 18887 18196 18896
rect 18144 18853 18153 18887
rect 18153 18853 18187 18887
rect 18187 18853 18196 18887
rect 18144 18844 18196 18853
rect 18328 18844 18380 18896
rect 18788 18844 18840 18896
rect 20260 18912 20312 18964
rect 21916 18955 21968 18964
rect 21916 18921 21925 18955
rect 21925 18921 21959 18955
rect 21959 18921 21968 18955
rect 21916 18912 21968 18921
rect 26056 18912 26108 18964
rect 20536 18844 20588 18896
rect 17776 18708 17828 18760
rect 19616 18708 19668 18760
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 23572 18776 23624 18828
rect 15016 18572 15068 18624
rect 18880 18640 18932 18692
rect 22192 18640 22244 18692
rect 22284 18640 22336 18692
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 17132 18572 17184 18624
rect 20168 18615 20220 18624
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20168 18572 20220 18581
rect 20904 18572 20956 18624
rect 22376 18572 22428 18624
rect 23572 18572 23624 18624
rect 24216 18572 24268 18624
rect 25504 18572 25556 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 9680 18368 9732 18420
rect 10324 18368 10376 18420
rect 10508 18368 10560 18420
rect 11520 18368 11572 18420
rect 4528 18343 4580 18352
rect 4528 18309 4537 18343
rect 4537 18309 4571 18343
rect 4571 18309 4580 18343
rect 4528 18300 4580 18309
rect 8392 18300 8444 18352
rect 8576 18300 8628 18352
rect 9956 18300 10008 18352
rect 12808 18300 12860 18352
rect 13452 18368 13504 18420
rect 14372 18368 14424 18420
rect 19248 18368 19300 18420
rect 19984 18368 20036 18420
rect 22100 18368 22152 18420
rect 13820 18300 13872 18352
rect 14832 18300 14884 18352
rect 17132 18343 17184 18352
rect 17132 18309 17141 18343
rect 17141 18309 17175 18343
rect 17175 18309 17184 18343
rect 17132 18300 17184 18309
rect 18420 18300 18472 18352
rect 18604 18300 18656 18352
rect 3792 18071 3844 18080
rect 3792 18037 3801 18071
rect 3801 18037 3835 18071
rect 3835 18037 3844 18071
rect 3792 18028 3844 18037
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 7288 18232 7340 18284
rect 11428 18232 11480 18284
rect 11888 18232 11940 18284
rect 12164 18232 12216 18284
rect 12072 18164 12124 18216
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 13452 18207 13504 18216
rect 13452 18173 13461 18207
rect 13461 18173 13495 18207
rect 13495 18173 13504 18207
rect 13452 18164 13504 18173
rect 15292 18232 15344 18284
rect 15476 18232 15528 18284
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 18880 18232 18932 18284
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 22376 18300 22428 18352
rect 23296 18232 23348 18284
rect 16028 18096 16080 18148
rect 25596 18164 25648 18216
rect 22008 18096 22060 18148
rect 23480 18096 23532 18148
rect 13912 18071 13964 18080
rect 13912 18037 13921 18071
rect 13921 18037 13955 18071
rect 13955 18037 13964 18071
rect 13912 18028 13964 18037
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 20168 18028 20220 18080
rect 22100 18028 22152 18080
rect 22836 18028 22888 18080
rect 25136 18028 25188 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 7840 17824 7892 17876
rect 9312 17824 9364 17876
rect 10968 17824 11020 17876
rect 11336 17824 11388 17876
rect 12164 17824 12216 17876
rect 12348 17824 12400 17876
rect 12808 17824 12860 17876
rect 13268 17824 13320 17876
rect 15200 17824 15252 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 20996 17824 21048 17876
rect 5448 17688 5500 17740
rect 5632 17620 5684 17672
rect 12440 17756 12492 17808
rect 6460 17731 6512 17740
rect 6460 17697 6469 17731
rect 6469 17697 6503 17731
rect 6503 17697 6512 17731
rect 6460 17688 6512 17697
rect 7748 17688 7800 17740
rect 9128 17688 9180 17740
rect 6552 17552 6604 17604
rect 7472 17620 7524 17672
rect 11336 17688 11388 17740
rect 14556 17756 14608 17808
rect 6828 17484 6880 17536
rect 6920 17484 6972 17536
rect 8484 17552 8536 17604
rect 9588 17595 9640 17604
rect 9588 17561 9597 17595
rect 9597 17561 9631 17595
rect 9631 17561 9640 17595
rect 9588 17552 9640 17561
rect 13268 17620 13320 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 15936 17688 15988 17740
rect 17592 17688 17644 17740
rect 18604 17731 18656 17740
rect 18604 17697 18613 17731
rect 18613 17697 18647 17731
rect 18647 17697 18656 17731
rect 18604 17688 18656 17697
rect 19064 17688 19116 17740
rect 23572 17688 23624 17740
rect 24860 17688 24912 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 15752 17620 15804 17672
rect 17776 17620 17828 17672
rect 18328 17620 18380 17672
rect 18696 17620 18748 17672
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 21456 17620 21508 17672
rect 22560 17620 22612 17672
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 9680 17484 9732 17536
rect 11244 17552 11296 17604
rect 11704 17484 11756 17536
rect 12072 17484 12124 17536
rect 13452 17595 13504 17604
rect 13452 17561 13461 17595
rect 13461 17561 13495 17595
rect 13495 17561 13504 17595
rect 13452 17552 13504 17561
rect 13912 17552 13964 17604
rect 16396 17552 16448 17604
rect 15476 17484 15528 17536
rect 16764 17527 16816 17536
rect 16764 17493 16773 17527
rect 16773 17493 16807 17527
rect 16807 17493 16816 17527
rect 16764 17484 16816 17493
rect 16948 17484 17000 17536
rect 17132 17484 17184 17536
rect 17316 17484 17368 17536
rect 17960 17484 18012 17536
rect 18328 17484 18380 17536
rect 19064 17484 19116 17536
rect 24584 17527 24636 17536
rect 24584 17493 24593 17527
rect 24593 17493 24627 17527
rect 24627 17493 24636 17527
rect 24584 17484 24636 17493
rect 24676 17484 24728 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 5356 17280 5408 17332
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 6276 17280 6328 17332
rect 8944 17280 8996 17332
rect 9956 17323 10008 17332
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 10048 17280 10100 17332
rect 12808 17280 12860 17332
rect 15568 17280 15620 17332
rect 15936 17280 15988 17332
rect 6828 17212 6880 17264
rect 9128 17212 9180 17264
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5908 17144 5960 17196
rect 8944 17144 8996 17196
rect 4436 17076 4488 17128
rect 5816 17076 5868 17128
rect 8300 17076 8352 17128
rect 9864 17212 9916 17264
rect 11336 17212 11388 17264
rect 11704 17212 11756 17264
rect 12532 17212 12584 17264
rect 9404 17076 9456 17128
rect 10324 17076 10376 17128
rect 11980 17144 12032 17196
rect 13912 17144 13964 17196
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 11520 17008 11572 17060
rect 2688 16940 2740 16992
rect 3608 16940 3660 16992
rect 6736 16940 6788 16992
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 8300 16940 8352 16992
rect 9680 16940 9732 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 12624 17076 12676 17128
rect 14372 17076 14424 17128
rect 14740 17076 14792 17128
rect 11888 17008 11940 17060
rect 17776 17144 17828 17196
rect 17500 17119 17552 17128
rect 17500 17085 17509 17119
rect 17509 17085 17543 17119
rect 17543 17085 17552 17119
rect 17500 17076 17552 17085
rect 17868 17076 17920 17128
rect 22192 17212 22244 17264
rect 22928 17323 22980 17332
rect 22928 17289 22937 17323
rect 22937 17289 22971 17323
rect 22971 17289 22980 17323
rect 22928 17280 22980 17289
rect 23848 17280 23900 17332
rect 24308 17212 24360 17264
rect 21272 17144 21324 17196
rect 21456 17187 21508 17196
rect 21456 17153 21465 17187
rect 21465 17153 21499 17187
rect 21499 17153 21508 17187
rect 21456 17144 21508 17153
rect 22008 17144 22060 17196
rect 23388 17144 23440 17196
rect 24032 17144 24084 17196
rect 23480 17076 23532 17128
rect 25136 17144 25188 17196
rect 24768 17119 24820 17128
rect 24768 17085 24777 17119
rect 24777 17085 24811 17119
rect 24811 17085 24820 17119
rect 24768 17076 24820 17085
rect 18420 17008 18472 17060
rect 22468 17051 22520 17060
rect 22468 17017 22477 17051
rect 22477 17017 22511 17051
rect 22511 17017 22520 17051
rect 22468 17008 22520 17017
rect 14648 16940 14700 16992
rect 14740 16940 14792 16992
rect 16948 16940 17000 16992
rect 17408 16940 17460 16992
rect 17500 16940 17552 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 5632 16736 5684 16788
rect 5540 16668 5592 16720
rect 6000 16668 6052 16720
rect 7748 16736 7800 16788
rect 4344 16600 4396 16652
rect 8300 16668 8352 16720
rect 6736 16600 6788 16652
rect 11060 16668 11112 16720
rect 13912 16736 13964 16788
rect 17224 16736 17276 16788
rect 19708 16736 19760 16788
rect 20812 16736 20864 16788
rect 22192 16779 22244 16788
rect 22192 16745 22201 16779
rect 22201 16745 22235 16779
rect 22235 16745 22244 16779
rect 22192 16736 22244 16745
rect 5908 16575 5960 16584
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 9220 16600 9272 16652
rect 9496 16532 9548 16584
rect 11152 16600 11204 16652
rect 12072 16668 12124 16720
rect 13360 16668 13412 16720
rect 14556 16668 14608 16720
rect 16028 16668 16080 16720
rect 11980 16532 12032 16584
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 14004 16600 14056 16652
rect 14188 16600 14240 16652
rect 16304 16600 16356 16652
rect 16856 16600 16908 16652
rect 18420 16600 18472 16652
rect 14280 16532 14332 16584
rect 6920 16464 6972 16516
rect 8576 16464 8628 16516
rect 9680 16464 9732 16516
rect 14832 16464 14884 16516
rect 15200 16464 15252 16516
rect 17224 16532 17276 16584
rect 18696 16600 18748 16652
rect 24676 16668 24728 16720
rect 20628 16600 20680 16652
rect 7932 16396 7984 16448
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 8852 16396 8904 16448
rect 10048 16396 10100 16448
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 11520 16396 11572 16448
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13360 16396 13412 16448
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 16672 16439 16724 16448
rect 16672 16405 16681 16439
rect 16681 16405 16715 16439
rect 16715 16405 16724 16439
rect 18880 16464 18932 16516
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 21548 16575 21600 16584
rect 21548 16541 21557 16575
rect 21557 16541 21591 16575
rect 21591 16541 21600 16575
rect 21548 16532 21600 16541
rect 16672 16396 16724 16405
rect 17132 16396 17184 16448
rect 20720 16396 20772 16448
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 21640 16396 21692 16448
rect 25964 16532 26016 16584
rect 25044 16464 25096 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 2044 16192 2096 16244
rect 4436 16192 4488 16244
rect 5540 16192 5592 16244
rect 6644 16192 6696 16244
rect 7748 16192 7800 16244
rect 9956 16192 10008 16244
rect 10692 16192 10744 16244
rect 3792 16124 3844 16176
rect 8116 16124 8168 16176
rect 8300 16124 8352 16176
rect 8484 16124 8536 16176
rect 10140 16124 10192 16176
rect 10784 16167 10836 16176
rect 10784 16133 10793 16167
rect 10793 16133 10827 16167
rect 10827 16133 10836 16167
rect 10784 16124 10836 16133
rect 11060 16124 11112 16176
rect 12256 16124 12308 16176
rect 13360 16124 13412 16176
rect 13544 16124 13596 16176
rect 14004 16124 14056 16176
rect 14832 16192 14884 16244
rect 16212 16192 16264 16244
rect 16488 16192 16540 16244
rect 21364 16192 21416 16244
rect 664 16056 716 16108
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 6184 16056 6236 16108
rect 7748 16056 7800 16108
rect 848 15988 900 16040
rect 6368 15988 6420 16040
rect 6644 15988 6696 16040
rect 7288 15988 7340 16040
rect 11520 16056 11572 16108
rect 2504 15920 2556 15972
rect 7840 15920 7892 15972
rect 7932 15920 7984 15972
rect 9772 15988 9824 16040
rect 2136 15852 2188 15904
rect 4160 15852 4212 15904
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 6920 15852 6972 15904
rect 8392 15852 8444 15904
rect 10140 15852 10192 15904
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 13084 15920 13136 15972
rect 13820 15920 13872 15972
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 15016 16124 15068 16176
rect 15200 16124 15252 16176
rect 18236 16124 18288 16176
rect 18788 16124 18840 16176
rect 20812 16124 20864 16176
rect 16396 16056 16448 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 25136 16167 25188 16176
rect 25136 16133 25145 16167
rect 25145 16133 25179 16167
rect 25179 16133 25188 16167
rect 25136 16124 25188 16133
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 15292 15963 15344 15972
rect 15292 15929 15301 15963
rect 15301 15929 15335 15963
rect 15335 15929 15344 15963
rect 15292 15920 15344 15929
rect 15752 16031 15804 16040
rect 15752 15997 15761 16031
rect 15761 15997 15795 16031
rect 15795 15997 15804 16031
rect 15752 15988 15804 15997
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 19340 15988 19392 16040
rect 15936 15920 15988 15972
rect 16212 15920 16264 15972
rect 11980 15852 12032 15904
rect 12716 15852 12768 15904
rect 13728 15852 13780 15904
rect 15016 15895 15068 15904
rect 15016 15861 15025 15895
rect 15025 15861 15059 15895
rect 15059 15861 15068 15895
rect 15016 15852 15068 15861
rect 16856 15852 16908 15904
rect 18420 15920 18472 15972
rect 21272 15988 21324 16040
rect 21640 15988 21692 16040
rect 23296 16031 23348 16040
rect 23296 15997 23305 16031
rect 23305 15997 23339 16031
rect 23339 15997 23348 16031
rect 23296 15988 23348 15997
rect 21824 15920 21876 15972
rect 20444 15852 20496 15904
rect 20812 15852 20864 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 572 15648 624 15700
rect 5356 15648 5408 15700
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 3424 15580 3476 15632
rect 3332 15512 3384 15564
rect 756 15444 808 15496
rect 4436 15487 4488 15496
rect 4436 15453 4445 15487
rect 4445 15453 4479 15487
rect 4479 15453 4488 15487
rect 4436 15444 4488 15453
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9036 15648 9088 15700
rect 9496 15648 9548 15700
rect 9404 15580 9456 15632
rect 6644 15555 6696 15564
rect 6644 15521 6653 15555
rect 6653 15521 6687 15555
rect 6687 15521 6696 15555
rect 6644 15512 6696 15521
rect 7288 15512 7340 15564
rect 11612 15648 11664 15700
rect 12256 15648 12308 15700
rect 16212 15648 16264 15700
rect 10140 15580 10192 15632
rect 8576 15444 8628 15496
rect 8760 15444 8812 15496
rect 11152 15512 11204 15564
rect 1032 15376 1084 15428
rect 3976 15376 4028 15428
rect 4252 15376 4304 15428
rect 7012 15376 7064 15428
rect 8484 15376 8536 15428
rect 9496 15376 9548 15428
rect 11060 15376 11112 15428
rect 12072 15512 12124 15564
rect 13268 15512 13320 15564
rect 12164 15444 12216 15496
rect 13176 15444 13228 15496
rect 13636 15555 13688 15564
rect 13636 15521 13645 15555
rect 13645 15521 13679 15555
rect 13679 15521 13688 15555
rect 13636 15512 13688 15521
rect 13728 15512 13780 15564
rect 16304 15555 16356 15564
rect 16304 15521 16313 15555
rect 16313 15521 16347 15555
rect 16347 15521 16356 15555
rect 16304 15512 16356 15521
rect 19064 15512 19116 15564
rect 20628 15512 20680 15564
rect 21824 15512 21876 15564
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 19248 15444 19300 15496
rect 25228 15444 25280 15496
rect 480 15308 532 15360
rect 2044 15351 2096 15360
rect 2044 15317 2053 15351
rect 2053 15317 2087 15351
rect 2087 15317 2096 15351
rect 2044 15308 2096 15317
rect 2228 15351 2280 15360
rect 2228 15317 2237 15351
rect 2237 15317 2271 15351
rect 2271 15317 2280 15351
rect 2228 15308 2280 15317
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 2872 15308 2924 15360
rect 3700 15308 3752 15360
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 7104 15308 7156 15360
rect 10140 15308 10192 15360
rect 10968 15308 11020 15360
rect 12164 15351 12216 15360
rect 12164 15317 12173 15351
rect 12173 15317 12207 15351
rect 12207 15317 12216 15351
rect 12164 15308 12216 15317
rect 12532 15308 12584 15360
rect 15936 15376 15988 15428
rect 18236 15376 18288 15428
rect 18788 15419 18840 15428
rect 18788 15385 18797 15419
rect 18797 15385 18831 15419
rect 18831 15385 18840 15419
rect 18788 15376 18840 15385
rect 19524 15419 19576 15428
rect 19524 15385 19533 15419
rect 19533 15385 19567 15419
rect 19567 15385 19576 15419
rect 19524 15376 19576 15385
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 19892 15376 19944 15428
rect 25044 15376 25096 15428
rect 13636 15308 13688 15360
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 15016 15308 15068 15360
rect 16028 15308 16080 15360
rect 16856 15308 16908 15360
rect 17592 15308 17644 15360
rect 20076 15308 20128 15360
rect 20996 15308 21048 15360
rect 25228 15308 25280 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 4436 15104 4488 15156
rect 5448 15104 5500 15156
rect 8944 15104 8996 15156
rect 9312 15104 9364 15156
rect 9588 15104 9640 15156
rect 14464 15104 14516 15156
rect 15568 15104 15620 15156
rect 16396 15104 16448 15156
rect 18328 15104 18380 15156
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 3884 14968 3936 15020
rect 8392 15036 8444 15088
rect 8576 15036 8628 15088
rect 9956 15036 10008 15088
rect 10324 15036 10376 15088
rect 11060 15036 11112 15088
rect 6000 14968 6052 15020
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7840 14968 7892 15020
rect 9588 14968 9640 15020
rect 11428 14968 11480 15020
rect 12716 14968 12768 15020
rect 1216 14900 1268 14952
rect 4344 14900 4396 14952
rect 5448 14900 5500 14952
rect 940 14832 992 14884
rect 8944 14900 8996 14952
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 15292 14968 15344 15020
rect 16580 14968 16632 15020
rect 6092 14832 6144 14884
rect 6552 14832 6604 14884
rect 6828 14832 6880 14884
rect 7748 14832 7800 14884
rect 13912 14900 13964 14952
rect 14188 14900 14240 14952
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 15016 14900 15068 14952
rect 16212 14900 16264 14952
rect 18604 14968 18656 15020
rect 20628 15104 20680 15156
rect 20996 15104 21048 15156
rect 20076 15036 20128 15088
rect 20904 15036 20956 15088
rect 24032 15147 24084 15156
rect 24032 15113 24041 15147
rect 24041 15113 24075 15147
rect 24075 15113 24084 15147
rect 24032 15104 24084 15113
rect 22376 15036 22428 15088
rect 24400 15011 24452 15020
rect 24400 14977 24409 15011
rect 24409 14977 24443 15011
rect 24443 14977 24452 15011
rect 24400 14968 24452 14977
rect 24676 15011 24728 15020
rect 24676 14977 24685 15011
rect 24685 14977 24719 15011
rect 24719 14977 24728 15011
rect 24676 14968 24728 14977
rect 17684 14900 17736 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 1952 14764 2004 14816
rect 2044 14764 2096 14816
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 3424 14764 3476 14816
rect 6276 14764 6328 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 8760 14764 8812 14816
rect 11796 14764 11848 14816
rect 15844 14832 15896 14884
rect 16120 14832 16172 14884
rect 20628 14900 20680 14952
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 20720 14832 20772 14884
rect 20904 14832 20956 14884
rect 13360 14764 13412 14816
rect 13452 14764 13504 14816
rect 13636 14764 13688 14816
rect 14740 14764 14792 14816
rect 18236 14764 18288 14816
rect 20628 14764 20680 14816
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 21640 14764 21692 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 4068 14560 4120 14612
rect 7012 14560 7064 14612
rect 7564 14560 7616 14612
rect 12624 14603 12676 14612
rect 12624 14569 12633 14603
rect 12633 14569 12667 14603
rect 12667 14569 12676 14603
rect 12624 14560 12676 14569
rect 13176 14560 13228 14612
rect 15568 14560 15620 14612
rect 16580 14603 16632 14612
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 22560 14560 22612 14612
rect 23664 14560 23716 14612
rect 2320 14492 2372 14544
rect 4436 14492 4488 14544
rect 5172 14492 5224 14544
rect 6000 14492 6052 14544
rect 7380 14492 7432 14544
rect 9588 14492 9640 14544
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 2688 14356 2740 14408
rect 6920 14424 6972 14476
rect 3884 14356 3936 14408
rect 8944 14424 8996 14476
rect 9312 14424 9364 14476
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 11704 14424 11756 14476
rect 11980 14424 12032 14476
rect 13636 14492 13688 14544
rect 14004 14492 14056 14544
rect 14188 14535 14240 14544
rect 14188 14501 14197 14535
rect 14197 14501 14231 14535
rect 14231 14501 14240 14535
rect 14188 14492 14240 14501
rect 14648 14492 14700 14544
rect 15752 14492 15804 14544
rect 13912 14467 13964 14476
rect 13912 14433 13921 14467
rect 13921 14433 13955 14467
rect 13955 14433 13964 14467
rect 13912 14424 13964 14433
rect 4068 14288 4120 14340
rect 1400 14220 1452 14272
rect 1860 14263 1912 14272
rect 1860 14229 1869 14263
rect 1869 14229 1903 14263
rect 1903 14229 1912 14263
rect 1860 14220 1912 14229
rect 5264 14331 5316 14340
rect 5264 14297 5273 14331
rect 5273 14297 5307 14331
rect 5307 14297 5316 14331
rect 5264 14288 5316 14297
rect 7104 14288 7156 14340
rect 7380 14288 7432 14340
rect 7656 14288 7708 14340
rect 9772 14356 9824 14408
rect 12716 14356 12768 14408
rect 14188 14356 14240 14408
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 15568 14424 15620 14476
rect 21732 14492 21784 14544
rect 16672 14424 16724 14476
rect 17776 14424 17828 14476
rect 20076 14467 20128 14476
rect 20076 14433 20085 14467
rect 20085 14433 20119 14467
rect 20119 14433 20128 14467
rect 20076 14424 20128 14433
rect 21640 14467 21692 14476
rect 21640 14433 21649 14467
rect 21649 14433 21683 14467
rect 21683 14433 21692 14467
rect 21640 14424 21692 14433
rect 22008 14424 22060 14476
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16856 14356 16908 14408
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 19524 14399 19576 14408
rect 19524 14365 19533 14399
rect 19533 14365 19567 14399
rect 19567 14365 19576 14399
rect 19524 14356 19576 14365
rect 20904 14356 20956 14408
rect 25136 14356 25188 14408
rect 6552 14220 6604 14272
rect 6736 14220 6788 14272
rect 7748 14220 7800 14272
rect 9772 14220 9824 14272
rect 10508 14220 10560 14272
rect 12072 14288 12124 14340
rect 12532 14288 12584 14340
rect 13912 14288 13964 14340
rect 14832 14288 14884 14340
rect 16028 14288 16080 14340
rect 17500 14288 17552 14340
rect 11980 14220 12032 14272
rect 13452 14220 13504 14272
rect 14280 14220 14332 14272
rect 15476 14220 15528 14272
rect 16212 14220 16264 14272
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 17684 14220 17736 14229
rect 18420 14220 18472 14272
rect 20904 14220 20956 14272
rect 22008 14288 22060 14340
rect 23020 14288 23072 14340
rect 22192 14220 22244 14272
rect 25044 14220 25096 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 1768 14016 1820 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6552 14016 6604 14068
rect 5724 13948 5776 14000
rect 2780 13880 2832 13932
rect 3884 13880 3936 13932
rect 4252 13923 4304 13932
rect 4252 13889 4261 13923
rect 4261 13889 4295 13923
rect 4295 13889 4304 13923
rect 4252 13880 4304 13889
rect 6276 13880 6328 13932
rect 9404 14016 9456 14068
rect 9496 14016 9548 14068
rect 10048 14016 10100 14068
rect 10876 14059 10928 14068
rect 7748 13948 7800 14000
rect 2136 13812 2188 13864
rect 10232 13948 10284 14000
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 13360 14016 13412 14068
rect 15200 14016 15252 14068
rect 17500 14016 17552 14068
rect 18512 14016 18564 14068
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 19340 14059 19392 14068
rect 19340 14025 19349 14059
rect 19349 14025 19383 14059
rect 19383 14025 19392 14059
rect 19340 14016 19392 14025
rect 19432 14016 19484 14068
rect 23940 14016 23992 14068
rect 25780 14016 25832 14068
rect 10692 13880 10744 13932
rect 8392 13812 8444 13864
rect 9128 13812 9180 13864
rect 8024 13744 8076 13796
rect 8760 13744 8812 13796
rect 9588 13744 9640 13796
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 11796 13880 11848 13932
rect 14280 13991 14332 14000
rect 14280 13957 14289 13991
rect 14289 13957 14323 13991
rect 14323 13957 14332 13991
rect 14280 13948 14332 13957
rect 14832 13948 14884 14000
rect 8392 13676 8444 13728
rect 8576 13676 8628 13728
rect 10232 13744 10284 13796
rect 10692 13744 10744 13796
rect 10784 13744 10836 13796
rect 11428 13812 11480 13864
rect 11980 13812 12032 13864
rect 13452 13880 13504 13932
rect 12256 13744 12308 13796
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 14648 13812 14700 13864
rect 19524 13948 19576 14000
rect 22100 13991 22152 14000
rect 22100 13957 22109 13991
rect 22109 13957 22143 13991
rect 22143 13957 22152 13991
rect 22100 13948 22152 13957
rect 16396 13923 16448 13932
rect 15384 13744 15436 13796
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 16396 13880 16448 13889
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 17868 13880 17920 13932
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 18972 13880 19024 13932
rect 20444 13880 20496 13932
rect 21824 13880 21876 13932
rect 23020 13948 23072 14000
rect 23848 13948 23900 14000
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 16028 13812 16080 13821
rect 15936 13744 15988 13796
rect 9956 13676 10008 13728
rect 13360 13676 13412 13728
rect 13452 13676 13504 13728
rect 16028 13676 16080 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16580 13676 16632 13728
rect 17592 13744 17644 13796
rect 20628 13812 20680 13864
rect 20904 13855 20956 13864
rect 20904 13821 20913 13855
rect 20913 13821 20947 13855
rect 20947 13821 20956 13855
rect 20904 13812 20956 13821
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 24492 13812 24544 13864
rect 21732 13744 21784 13796
rect 25228 13744 25280 13796
rect 25412 13744 25464 13796
rect 21272 13676 21324 13728
rect 24860 13676 24912 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 2596 13472 2648 13524
rect 5632 13404 5684 13456
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 7748 13472 7800 13524
rect 7932 13472 7984 13524
rect 9220 13472 9272 13524
rect 9864 13472 9916 13524
rect 10508 13472 10560 13524
rect 12256 13472 12308 13524
rect 5540 13336 5592 13388
rect 5908 13336 5960 13388
rect 11980 13404 12032 13456
rect 12440 13472 12492 13524
rect 13728 13472 13780 13524
rect 14096 13472 14148 13524
rect 16028 13472 16080 13524
rect 18880 13515 18932 13524
rect 18880 13481 18889 13515
rect 18889 13481 18923 13515
rect 18923 13481 18932 13515
rect 18880 13472 18932 13481
rect 19340 13515 19392 13524
rect 19340 13481 19349 13515
rect 19349 13481 19383 13515
rect 19383 13481 19392 13515
rect 19340 13472 19392 13481
rect 21088 13472 21140 13524
rect 22652 13472 22704 13524
rect 24124 13472 24176 13524
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 4160 13268 4212 13320
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 4528 13311 4580 13320
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 3424 13200 3476 13252
rect 5172 13243 5224 13252
rect 5172 13209 5181 13243
rect 5181 13209 5215 13243
rect 5215 13209 5224 13243
rect 5172 13200 5224 13209
rect 5448 13200 5500 13252
rect 8024 13268 8076 13320
rect 8116 13268 8168 13320
rect 9312 13336 9364 13388
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 9772 13336 9824 13388
rect 12072 13336 12124 13388
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 12348 13379 12400 13388
rect 12348 13345 12357 13379
rect 12357 13345 12391 13379
rect 12391 13345 12400 13379
rect 12348 13336 12400 13345
rect 8944 13268 8996 13320
rect 9128 13268 9180 13320
rect 12440 13268 12492 13320
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 17040 13404 17092 13456
rect 18512 13404 18564 13456
rect 16028 13336 16080 13388
rect 16120 13336 16172 13388
rect 19432 13336 19484 13388
rect 19524 13336 19576 13388
rect 20628 13336 20680 13388
rect 15936 13268 15988 13320
rect 17684 13268 17736 13320
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 7472 13200 7524 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 3884 13132 3936 13184
rect 5356 13132 5408 13184
rect 7748 13132 7800 13184
rect 8760 13200 8812 13252
rect 7932 13132 7984 13184
rect 8944 13132 8996 13184
rect 9772 13132 9824 13184
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 12072 13200 12124 13252
rect 11980 13132 12032 13184
rect 12900 13132 12952 13184
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 14096 13200 14148 13252
rect 15476 13200 15528 13252
rect 19248 13268 19300 13320
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21364 13200 21416 13252
rect 21916 13268 21968 13320
rect 23940 13336 23992 13388
rect 23756 13268 23808 13320
rect 24216 13268 24268 13320
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 24492 13200 24544 13252
rect 15108 13132 15160 13184
rect 15200 13132 15252 13184
rect 15384 13132 15436 13184
rect 15568 13132 15620 13184
rect 16856 13132 16908 13184
rect 17868 13132 17920 13184
rect 19064 13132 19116 13184
rect 19340 13132 19392 13184
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 22560 13132 22612 13184
rect 22928 13132 22980 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 1124 12588 1176 12640
rect 3608 12928 3660 12980
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 4804 12928 4856 12980
rect 7748 12928 7800 12980
rect 8668 12928 8720 12980
rect 9404 12928 9456 12980
rect 10508 12928 10560 12980
rect 12164 12928 12216 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 14188 12928 14240 12980
rect 16580 12928 16632 12980
rect 9772 12860 9824 12912
rect 10140 12860 10192 12912
rect 11888 12860 11940 12912
rect 12348 12860 12400 12912
rect 14372 12860 14424 12912
rect 3792 12792 3844 12844
rect 5080 12792 5132 12844
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8576 12792 8628 12844
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 11980 12792 12032 12844
rect 8484 12724 8536 12776
rect 1768 12656 1820 12708
rect 5448 12656 5500 12708
rect 5632 12656 5684 12708
rect 3792 12631 3844 12640
rect 3792 12597 3801 12631
rect 3801 12597 3835 12631
rect 3835 12597 3844 12631
rect 3792 12588 3844 12597
rect 5356 12588 5408 12640
rect 6000 12631 6052 12640
rect 6000 12597 6009 12631
rect 6009 12597 6043 12631
rect 6043 12597 6052 12631
rect 6000 12588 6052 12597
rect 6368 12588 6420 12640
rect 6552 12588 6604 12640
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 7748 12588 7800 12640
rect 8208 12656 8260 12708
rect 8760 12656 8812 12708
rect 11704 12656 11756 12708
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 18144 12928 18196 12980
rect 18420 12928 18472 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 19432 12928 19484 12980
rect 20628 12928 20680 12980
rect 21916 12928 21968 12980
rect 17868 12860 17920 12912
rect 18880 12860 18932 12912
rect 19064 12903 19116 12912
rect 19064 12869 19073 12903
rect 19073 12869 19107 12903
rect 19107 12869 19116 12903
rect 19064 12860 19116 12869
rect 19340 12860 19392 12912
rect 19616 12903 19668 12912
rect 19616 12869 19625 12903
rect 19625 12869 19659 12903
rect 19659 12869 19668 12903
rect 19616 12860 19668 12869
rect 19800 12860 19852 12912
rect 22008 12860 22060 12912
rect 22376 12860 22428 12912
rect 23296 12903 23348 12912
rect 23296 12869 23305 12903
rect 23305 12869 23339 12903
rect 23339 12869 23348 12903
rect 23296 12860 23348 12869
rect 23848 12860 23900 12912
rect 24584 12860 24636 12912
rect 16212 12792 16264 12844
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16120 12724 16172 12733
rect 12164 12656 12216 12708
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 11612 12588 11664 12640
rect 14188 12588 14240 12640
rect 14648 12588 14700 12640
rect 15108 12588 15160 12640
rect 16580 12588 16632 12640
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 17224 12724 17276 12776
rect 20444 12767 20496 12776
rect 20444 12733 20453 12767
rect 20453 12733 20487 12767
rect 20487 12733 20496 12767
rect 20444 12724 20496 12733
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 24860 12792 24912 12844
rect 21824 12724 21876 12776
rect 21916 12724 21968 12776
rect 22652 12724 22704 12776
rect 22836 12724 22888 12776
rect 23848 12724 23900 12776
rect 24492 12724 24544 12776
rect 18144 12656 18196 12708
rect 18512 12588 18564 12640
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 20720 12588 20772 12640
rect 21272 12588 21324 12640
rect 21456 12588 21508 12640
rect 21640 12588 21692 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 4528 12384 4580 12436
rect 7104 12384 7156 12436
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 4068 12248 4120 12300
rect 4712 12316 4764 12368
rect 9864 12384 9916 12436
rect 10600 12384 10652 12436
rect 11060 12384 11112 12436
rect 11520 12384 11572 12436
rect 13176 12384 13228 12436
rect 13820 12384 13872 12436
rect 14648 12384 14700 12436
rect 14832 12384 14884 12436
rect 14924 12384 14976 12436
rect 17224 12384 17276 12436
rect 17684 12384 17736 12436
rect 7748 12316 7800 12368
rect 10048 12316 10100 12368
rect 10784 12316 10836 12368
rect 11152 12316 11204 12368
rect 13636 12316 13688 12368
rect 18696 12384 18748 12436
rect 19800 12384 19852 12436
rect 4252 12180 4304 12232
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 6000 12180 6052 12232
rect 11244 12248 11296 12300
rect 8024 12180 8076 12232
rect 8208 12112 8260 12164
rect 8852 12180 8904 12232
rect 9772 12180 9824 12232
rect 11796 12248 11848 12300
rect 11980 12248 12032 12300
rect 12348 12248 12400 12300
rect 15016 12291 15068 12300
rect 15016 12257 15025 12291
rect 15025 12257 15059 12291
rect 15059 12257 15068 12291
rect 15016 12248 15068 12257
rect 15568 12248 15620 12300
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 3792 12044 3844 12096
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4712 12044 4764 12096
rect 8024 12044 8076 12096
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 8760 12044 8812 12096
rect 9680 12155 9732 12164
rect 9680 12121 9689 12155
rect 9689 12121 9723 12155
rect 9723 12121 9732 12155
rect 9680 12112 9732 12121
rect 10600 12155 10652 12164
rect 10600 12121 10609 12155
rect 10609 12121 10643 12155
rect 10643 12121 10652 12155
rect 10600 12112 10652 12121
rect 10692 12112 10744 12164
rect 12256 12180 12308 12232
rect 13452 12180 13504 12232
rect 14740 12180 14792 12232
rect 15108 12180 15160 12232
rect 11888 12112 11940 12164
rect 13728 12112 13780 12164
rect 14004 12112 14056 12164
rect 14648 12112 14700 12164
rect 16948 12180 17000 12232
rect 20260 12316 20312 12368
rect 18696 12248 18748 12300
rect 20904 12384 20956 12436
rect 22744 12384 22796 12436
rect 25320 12384 25372 12436
rect 22468 12316 22520 12368
rect 23480 12316 23532 12368
rect 20444 12291 20496 12300
rect 20444 12257 20453 12291
rect 20453 12257 20487 12291
rect 20487 12257 20496 12291
rect 20444 12248 20496 12257
rect 22652 12248 22704 12300
rect 24216 12248 24268 12300
rect 19524 12180 19576 12232
rect 12256 12044 12308 12096
rect 12348 12044 12400 12096
rect 13452 12044 13504 12096
rect 14188 12044 14240 12096
rect 15016 12044 15068 12096
rect 15384 12044 15436 12096
rect 19984 12112 20036 12164
rect 20168 12180 20220 12232
rect 20352 12180 20404 12232
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 25044 12180 25096 12232
rect 22008 12112 22060 12164
rect 17316 12044 17368 12096
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 18420 12044 18472 12096
rect 19432 12087 19484 12096
rect 19432 12053 19441 12087
rect 19441 12053 19475 12087
rect 19475 12053 19484 12087
rect 19432 12044 19484 12053
rect 20260 12044 20312 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 4804 11840 4856 11892
rect 5080 11883 5132 11892
rect 5080 11849 5089 11883
rect 5089 11849 5123 11883
rect 5123 11849 5132 11883
rect 5080 11840 5132 11849
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 3884 11704 3936 11756
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 9220 11840 9272 11892
rect 9588 11840 9640 11892
rect 10048 11840 10100 11892
rect 10692 11840 10744 11892
rect 10876 11840 10928 11892
rect 11152 11840 11204 11892
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 11888 11840 11940 11892
rect 12532 11840 12584 11892
rect 12624 11840 12676 11892
rect 13544 11840 13596 11892
rect 14280 11840 14332 11892
rect 14556 11840 14608 11892
rect 14648 11840 14700 11892
rect 15568 11840 15620 11892
rect 16028 11840 16080 11892
rect 6644 11772 6696 11824
rect 6828 11772 6880 11824
rect 8116 11772 8168 11824
rect 11428 11772 11480 11824
rect 11612 11772 11664 11824
rect 13360 11772 13412 11824
rect 13452 11772 13504 11824
rect 17408 11840 17460 11892
rect 17500 11840 17552 11892
rect 19432 11772 19484 11824
rect 20168 11772 20220 11824
rect 20352 11772 20404 11824
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 21732 11772 21784 11824
rect 24860 11772 24912 11824
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 10508 11704 10560 11756
rect 11520 11704 11572 11756
rect 12624 11704 12676 11756
rect 13176 11704 13228 11756
rect 13544 11704 13596 11756
rect 14004 11704 14056 11756
rect 14372 11704 14424 11756
rect 5908 11636 5960 11688
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 2136 11500 2188 11552
rect 3516 11568 3568 11620
rect 4528 11568 4580 11620
rect 6920 11611 6972 11620
rect 6920 11577 6929 11611
rect 6929 11577 6963 11611
rect 6963 11577 6972 11611
rect 6920 11568 6972 11577
rect 4160 11500 4212 11552
rect 4252 11500 4304 11552
rect 7104 11500 7156 11552
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 8116 11636 8168 11688
rect 8668 11636 8720 11688
rect 9404 11636 9456 11688
rect 10876 11636 10928 11688
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 8944 11568 8996 11620
rect 9220 11568 9272 11620
rect 13636 11568 13688 11620
rect 14188 11636 14240 11688
rect 14832 11747 14884 11756
rect 14832 11713 14841 11747
rect 14841 11713 14875 11747
rect 14875 11713 14884 11747
rect 14832 11704 14884 11713
rect 16028 11704 16080 11756
rect 18604 11704 18656 11756
rect 20260 11704 20312 11756
rect 20812 11704 20864 11756
rect 20996 11704 21048 11756
rect 23756 11704 23808 11756
rect 15016 11568 15068 11620
rect 18328 11636 18380 11688
rect 18512 11636 18564 11688
rect 20628 11636 20680 11688
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 8760 11500 8812 11552
rect 10416 11500 10468 11552
rect 11980 11500 12032 11552
rect 16212 11500 16264 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 20260 11543 20312 11552
rect 20260 11509 20269 11543
rect 20269 11509 20303 11543
rect 20303 11509 20312 11543
rect 20260 11500 20312 11509
rect 20352 11500 20404 11552
rect 23572 11500 23624 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 3884 11296 3936 11348
rect 6552 11296 6604 11348
rect 7656 11296 7708 11348
rect 8392 11296 8444 11348
rect 9496 11296 9548 11348
rect 10968 11296 11020 11348
rect 11888 11296 11940 11348
rect 14372 11296 14424 11348
rect 14464 11296 14516 11348
rect 15016 11296 15068 11348
rect 17500 11296 17552 11348
rect 17684 11296 17736 11348
rect 17868 11339 17920 11348
rect 17868 11305 17877 11339
rect 17877 11305 17911 11339
rect 17911 11305 17920 11339
rect 17868 11296 17920 11305
rect 18972 11296 19024 11348
rect 19340 11339 19392 11348
rect 19340 11305 19349 11339
rect 19349 11305 19383 11339
rect 19383 11305 19392 11339
rect 19340 11296 19392 11305
rect 21088 11296 21140 11348
rect 22744 11296 22796 11348
rect 4712 11228 4764 11280
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 2688 11024 2740 11076
rect 4068 11092 4120 11144
rect 4344 11092 4396 11144
rect 11612 11228 11664 11280
rect 11704 11228 11756 11280
rect 7288 11160 7340 11212
rect 7380 11160 7432 11212
rect 8208 11160 8260 11212
rect 8484 11160 8536 11212
rect 10324 11160 10376 11212
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 10968 11160 11020 11212
rect 11796 11160 11848 11212
rect 12716 11228 12768 11280
rect 13084 11228 13136 11280
rect 16028 11228 16080 11280
rect 16120 11228 16172 11280
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 13544 11160 13596 11212
rect 14832 11160 14884 11212
rect 15292 11160 15344 11212
rect 16212 11160 16264 11212
rect 6644 11092 6696 11144
rect 3240 11067 3292 11076
rect 3240 11033 3249 11067
rect 3249 11033 3283 11067
rect 3283 11033 3292 11067
rect 3240 11024 3292 11033
rect 1860 10956 1912 11008
rect 2780 10956 2832 11008
rect 4804 11024 4856 11076
rect 8392 11092 8444 11144
rect 8576 11092 8628 11144
rect 8852 11024 8904 11076
rect 8944 11024 8996 11076
rect 9864 11092 9916 11144
rect 13176 11092 13228 11144
rect 13360 11092 13412 11144
rect 10508 11024 10560 11076
rect 4712 10999 4764 11008
rect 4712 10965 4721 10999
rect 4721 10965 4755 10999
rect 4755 10965 4764 10999
rect 4712 10956 4764 10965
rect 4896 10956 4948 11008
rect 6184 10956 6236 11008
rect 10416 10956 10468 11008
rect 10692 10956 10744 11008
rect 11152 10956 11204 11008
rect 12164 10956 12216 11008
rect 12532 10956 12584 11008
rect 13636 11024 13688 11076
rect 16304 11092 16356 11144
rect 16764 11092 16816 11144
rect 19800 11228 19852 11280
rect 18604 11160 18656 11212
rect 18696 11203 18748 11212
rect 18696 11169 18705 11203
rect 18705 11169 18739 11203
rect 18739 11169 18748 11203
rect 18696 11160 18748 11169
rect 18972 11160 19024 11212
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 20260 11160 20312 11212
rect 17776 11092 17828 11144
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 14556 11024 14608 11076
rect 14832 11024 14884 11076
rect 15108 10956 15160 11008
rect 15292 11024 15344 11076
rect 15476 11024 15528 11076
rect 17684 11024 17736 11076
rect 18972 11024 19024 11076
rect 18512 10999 18564 11008
rect 18512 10965 18521 10999
rect 18521 10965 18555 10999
rect 18555 10965 18564 10999
rect 18512 10956 18564 10965
rect 20352 11024 20404 11076
rect 21640 11024 21692 11076
rect 24860 11024 24912 11076
rect 20168 10956 20220 11008
rect 20260 10956 20312 11008
rect 22284 10956 22336 11008
rect 23664 10956 23716 11008
rect 24492 10956 24544 11008
rect 25044 10956 25096 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 1860 10752 1912 10804
rect 1400 10684 1452 10736
rect 5264 10752 5316 10804
rect 4712 10684 4764 10736
rect 6736 10752 6788 10804
rect 8852 10795 8904 10804
rect 8852 10761 8861 10795
rect 8861 10761 8895 10795
rect 8895 10761 8904 10795
rect 8852 10752 8904 10761
rect 7288 10727 7340 10736
rect 7288 10693 7297 10727
rect 7297 10693 7331 10727
rect 7331 10693 7340 10727
rect 7288 10684 7340 10693
rect 7472 10727 7524 10736
rect 7472 10693 7481 10727
rect 7481 10693 7515 10727
rect 7515 10693 7524 10727
rect 7472 10684 7524 10693
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 2688 10455 2740 10464
rect 2688 10421 2697 10455
rect 2697 10421 2731 10455
rect 2731 10421 2740 10455
rect 2688 10412 2740 10421
rect 5908 10616 5960 10668
rect 6184 10616 6236 10668
rect 6920 10616 6972 10668
rect 8024 10616 8076 10668
rect 10876 10752 10928 10804
rect 11152 10752 11204 10804
rect 15292 10752 15344 10804
rect 15752 10752 15804 10804
rect 9312 10684 9364 10736
rect 10140 10684 10192 10736
rect 12072 10727 12124 10736
rect 12072 10693 12081 10727
rect 12081 10693 12115 10727
rect 12115 10693 12124 10727
rect 12072 10684 12124 10693
rect 11060 10616 11112 10668
rect 14372 10684 14424 10736
rect 15016 10684 15068 10736
rect 16028 10752 16080 10804
rect 17868 10752 17920 10804
rect 21916 10752 21968 10804
rect 16212 10684 16264 10736
rect 16488 10684 16540 10736
rect 15476 10616 15528 10668
rect 16396 10616 16448 10668
rect 16764 10616 16816 10668
rect 17592 10616 17644 10668
rect 18420 10616 18472 10668
rect 6000 10548 6052 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 4988 10480 5040 10532
rect 6736 10480 6788 10532
rect 11152 10548 11204 10600
rect 10876 10480 10928 10532
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 13360 10548 13412 10600
rect 13820 10548 13872 10600
rect 14280 10548 14332 10600
rect 14556 10591 14608 10600
rect 14556 10557 14565 10591
rect 14565 10557 14599 10591
rect 14599 10557 14608 10591
rect 14556 10548 14608 10557
rect 13544 10480 13596 10532
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 17316 10548 17368 10600
rect 19340 10616 19392 10668
rect 19156 10548 19208 10600
rect 16488 10480 16540 10532
rect 5080 10412 5132 10464
rect 5724 10412 5776 10464
rect 6920 10412 6972 10464
rect 7748 10412 7800 10464
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 8024 10412 8076 10464
rect 10232 10412 10284 10464
rect 10324 10412 10376 10464
rect 11796 10412 11848 10464
rect 11888 10412 11940 10464
rect 13176 10412 13228 10464
rect 13820 10412 13872 10464
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 14280 10412 14332 10464
rect 14832 10412 14884 10464
rect 14924 10412 14976 10464
rect 15108 10412 15160 10464
rect 18512 10480 18564 10532
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 20260 10727 20312 10736
rect 20260 10693 20269 10727
rect 20269 10693 20303 10727
rect 20303 10693 20312 10727
rect 20260 10684 20312 10693
rect 22376 10727 22428 10736
rect 22376 10693 22385 10727
rect 22385 10693 22419 10727
rect 22419 10693 22428 10727
rect 22376 10684 22428 10693
rect 23296 10727 23348 10736
rect 23296 10693 23305 10727
rect 23305 10693 23339 10727
rect 23339 10693 23348 10727
rect 23296 10684 23348 10693
rect 25044 10727 25096 10736
rect 25044 10693 25053 10727
rect 25053 10693 25087 10727
rect 25087 10693 25096 10727
rect 25044 10684 25096 10693
rect 20352 10616 20404 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 22560 10616 22612 10668
rect 22652 10616 22704 10668
rect 24400 10616 24452 10668
rect 19708 10480 19760 10532
rect 22284 10548 22336 10600
rect 22376 10480 22428 10532
rect 23480 10412 23532 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 5908 10208 5960 10260
rect 6000 10208 6052 10260
rect 1400 10072 1452 10124
rect 4252 10140 4304 10192
rect 7748 10140 7800 10192
rect 8392 10208 8444 10260
rect 8668 10208 8720 10260
rect 9128 10208 9180 10260
rect 1400 9936 1452 9988
rect 3424 10004 3476 10056
rect 3240 9979 3292 9988
rect 3240 9945 3249 9979
rect 3249 9945 3283 9979
rect 3283 9945 3292 9979
rect 3240 9936 3292 9945
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 5908 10004 5960 10056
rect 8484 10072 8536 10124
rect 9404 10072 9456 10124
rect 9772 10072 9824 10124
rect 7288 10004 7340 10056
rect 9036 10004 9088 10056
rect 10692 10208 10744 10260
rect 11520 10208 11572 10260
rect 12164 10208 12216 10260
rect 11152 10140 11204 10192
rect 12532 10140 12584 10192
rect 12716 10140 12768 10192
rect 14280 10208 14332 10260
rect 10876 10115 10928 10124
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 11244 10072 11296 10124
rect 11520 10072 11572 10124
rect 11612 10072 11664 10124
rect 14188 10140 14240 10192
rect 14372 10140 14424 10192
rect 15844 10208 15896 10260
rect 17132 10208 17184 10260
rect 17868 10208 17920 10260
rect 19708 10208 19760 10260
rect 19984 10208 20036 10260
rect 20720 10208 20772 10260
rect 20904 10208 20956 10260
rect 25688 10208 25740 10260
rect 16856 10140 16908 10192
rect 18696 10140 18748 10192
rect 22376 10183 22428 10192
rect 22376 10149 22385 10183
rect 22385 10149 22419 10183
rect 22419 10149 22428 10183
rect 22376 10140 22428 10149
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 4988 9868 5040 9920
rect 5448 9868 5500 9920
rect 7104 9936 7156 9988
rect 9496 9936 9548 9988
rect 7196 9868 7248 9920
rect 9588 9868 9640 9920
rect 10140 9936 10192 9988
rect 10784 9936 10836 9988
rect 13544 9936 13596 9988
rect 13820 10004 13872 10056
rect 16764 10004 16816 10056
rect 19248 10072 19300 10124
rect 23480 10115 23532 10124
rect 23480 10081 23489 10115
rect 23489 10081 23523 10115
rect 23523 10081 23532 10115
rect 23480 10072 23532 10081
rect 17684 10004 17736 10056
rect 18328 10004 18380 10056
rect 20628 10047 20680 10056
rect 20628 10013 20637 10047
rect 20637 10013 20671 10047
rect 20671 10013 20680 10047
rect 20628 10004 20680 10013
rect 22008 10004 22060 10056
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 24308 10004 24360 10056
rect 11060 9868 11112 9920
rect 11520 9868 11572 9920
rect 14740 9936 14792 9988
rect 16396 9936 16448 9988
rect 14556 9868 14608 9920
rect 14832 9868 14884 9920
rect 15660 9868 15712 9920
rect 16120 9868 16172 9920
rect 16764 9868 16816 9920
rect 17868 9868 17920 9920
rect 18328 9868 18380 9920
rect 18696 9868 18748 9920
rect 18972 9868 19024 9920
rect 19432 9868 19484 9920
rect 22284 9868 22336 9920
rect 22836 9868 22888 9920
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 1492 9528 1544 9580
rect 2228 9528 2280 9580
rect 3240 9639 3292 9648
rect 3240 9605 3249 9639
rect 3249 9605 3283 9639
rect 3283 9605 3292 9639
rect 3240 9596 3292 9605
rect 4436 9596 4488 9648
rect 4528 9596 4580 9648
rect 5264 9664 5316 9716
rect 8208 9664 8260 9716
rect 9036 9664 9088 9716
rect 10876 9664 10928 9716
rect 11244 9664 11296 9716
rect 12164 9664 12216 9716
rect 12256 9664 12308 9716
rect 6184 9596 6236 9648
rect 7288 9639 7340 9648
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 7656 9596 7708 9648
rect 9404 9596 9456 9648
rect 1860 9460 1912 9512
rect 4252 9528 4304 9580
rect 12440 9596 12492 9648
rect 14004 9664 14056 9716
rect 14648 9596 14700 9648
rect 7564 9460 7616 9512
rect 1308 9392 1360 9444
rect 2320 9392 2372 9444
rect 7380 9392 7432 9444
rect 10416 9528 10468 9580
rect 13452 9528 13504 9580
rect 8760 9460 8812 9512
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9772 9460 9824 9512
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 4068 9324 4120 9376
rect 4528 9324 4580 9376
rect 4988 9324 5040 9376
rect 7656 9324 7708 9376
rect 10140 9392 10192 9444
rect 10416 9392 10468 9444
rect 11612 9392 11664 9444
rect 11520 9324 11572 9376
rect 12624 9460 12676 9512
rect 13176 9460 13228 9512
rect 14372 9528 14424 9580
rect 15844 9596 15896 9648
rect 16212 9596 16264 9648
rect 16948 9639 17000 9648
rect 16948 9605 16957 9639
rect 16957 9605 16991 9639
rect 16991 9605 17000 9639
rect 16948 9596 17000 9605
rect 17224 9664 17276 9716
rect 20536 9664 20588 9716
rect 20720 9664 20772 9716
rect 24032 9664 24084 9716
rect 18420 9596 18472 9648
rect 19892 9596 19944 9648
rect 19984 9596 20036 9648
rect 14832 9460 14884 9512
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 12716 9324 12768 9376
rect 13728 9392 13780 9444
rect 14004 9392 14056 9444
rect 14188 9392 14240 9444
rect 14740 9392 14792 9444
rect 13452 9324 13504 9376
rect 16120 9392 16172 9444
rect 16304 9435 16356 9444
rect 16304 9401 16313 9435
rect 16313 9401 16347 9435
rect 16347 9401 16356 9435
rect 16304 9392 16356 9401
rect 16764 9392 16816 9444
rect 17592 9460 17644 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18328 9503 18380 9512
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 20352 9528 20404 9580
rect 19616 9460 19668 9512
rect 22744 9528 22796 9580
rect 23664 9528 23716 9580
rect 22284 9460 22336 9512
rect 23296 9503 23348 9512
rect 23296 9469 23305 9503
rect 23305 9469 23339 9503
rect 23339 9469 23348 9503
rect 23296 9460 23348 9469
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 20996 9392 21048 9444
rect 21548 9392 21600 9444
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17132 9324 17184 9376
rect 17500 9324 17552 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 18972 9324 19024 9376
rect 22468 9324 22520 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 4712 9120 4764 9172
rect 6644 9120 6696 9172
rect 8944 9120 8996 9172
rect 9128 9120 9180 9172
rect 12072 9120 12124 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 13636 9120 13688 9172
rect 15936 9163 15988 9172
rect 15936 9129 15945 9163
rect 15945 9129 15979 9163
rect 15979 9129 15988 9163
rect 15936 9120 15988 9129
rect 3516 9052 3568 9104
rect 4068 9052 4120 9104
rect 6368 9052 6420 9104
rect 10232 9052 10284 9104
rect 11796 9052 11848 9104
rect 12808 9052 12860 9104
rect 16028 9052 16080 9104
rect 2412 8984 2464 9036
rect 1676 8916 1728 8968
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 7196 8916 7248 8968
rect 1584 8848 1636 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 3148 8780 3200 8832
rect 6736 8848 6788 8900
rect 8852 8984 8904 9036
rect 8300 8916 8352 8968
rect 10600 8984 10652 9036
rect 11152 8984 11204 9036
rect 12348 8984 12400 9036
rect 12532 8984 12584 9036
rect 13820 8984 13872 9036
rect 14004 8984 14056 9036
rect 14188 8984 14240 9036
rect 14464 8984 14516 9036
rect 14924 8984 14976 9036
rect 15568 8984 15620 9036
rect 9496 8916 9548 8968
rect 10232 8848 10284 8900
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 12440 8916 12492 8968
rect 16120 8916 16172 8968
rect 11244 8848 11296 8900
rect 12256 8848 12308 8900
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 5356 8780 5408 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 9680 8780 9732 8832
rect 10784 8780 10836 8832
rect 13636 8780 13688 8832
rect 13728 8823 13780 8832
rect 13728 8789 13737 8823
rect 13737 8789 13771 8823
rect 13771 8789 13780 8823
rect 13728 8780 13780 8789
rect 14188 8848 14240 8900
rect 19800 9120 19852 9172
rect 19156 9052 19208 9104
rect 25228 9163 25280 9172
rect 25228 9129 25237 9163
rect 25237 9129 25271 9163
rect 25271 9129 25280 9163
rect 25228 9120 25280 9129
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 17408 9027 17460 9036
rect 17408 8993 17417 9027
rect 17417 8993 17451 9027
rect 17451 8993 17460 9027
rect 17408 8984 17460 8993
rect 17500 8984 17552 9036
rect 20628 8984 20680 9036
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 21916 8916 21968 8968
rect 22008 8916 22060 8968
rect 22652 8984 22704 9036
rect 24676 8916 24728 8968
rect 16488 8848 16540 8900
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 15200 8823 15252 8832
rect 15200 8789 15209 8823
rect 15209 8789 15243 8823
rect 15243 8789 15252 8823
rect 15200 8780 15252 8789
rect 16212 8780 16264 8832
rect 17500 8848 17552 8900
rect 17960 8848 18012 8900
rect 18696 8848 18748 8900
rect 16672 8780 16724 8832
rect 19248 8780 19300 8832
rect 19616 8780 19668 8832
rect 22100 8891 22152 8900
rect 22100 8857 22109 8891
rect 22109 8857 22143 8891
rect 22143 8857 22152 8891
rect 22100 8848 22152 8857
rect 22744 8780 22796 8832
rect 22836 8780 22888 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 3148 8576 3200 8628
rect 6828 8576 6880 8628
rect 7196 8619 7248 8628
rect 7196 8585 7205 8619
rect 7205 8585 7239 8619
rect 7239 8585 7248 8619
rect 7196 8576 7248 8585
rect 7472 8576 7524 8628
rect 7748 8576 7800 8628
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 1584 8440 1636 8492
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2780 8508 2832 8560
rect 3792 8508 3844 8560
rect 4160 8508 4212 8560
rect 5908 8508 5960 8560
rect 6368 8508 6420 8560
rect 6644 8508 6696 8560
rect 7564 8508 7616 8560
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 8576 8508 8628 8560
rect 13820 8576 13872 8628
rect 13912 8576 13964 8628
rect 14372 8619 14424 8628
rect 14372 8585 14381 8619
rect 14381 8585 14415 8619
rect 14415 8585 14424 8619
rect 14372 8576 14424 8585
rect 15108 8576 15160 8628
rect 16764 8576 16816 8628
rect 18328 8576 18380 8628
rect 20444 8576 20496 8628
rect 4068 8440 4120 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 2688 8347 2740 8356
rect 2688 8313 2697 8347
rect 2697 8313 2731 8347
rect 2731 8313 2740 8347
rect 2688 8304 2740 8313
rect 7472 8440 7524 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 10140 8440 10192 8492
rect 8392 8372 8444 8424
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 13636 8508 13688 8560
rect 14648 8508 14700 8560
rect 15568 8508 15620 8560
rect 16212 8508 16264 8560
rect 16948 8508 17000 8560
rect 17408 8508 17460 8560
rect 17500 8508 17552 8560
rect 19248 8508 19300 8560
rect 21548 8508 21600 8560
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 5356 8304 5408 8356
rect 1124 8236 1176 8288
rect 3884 8236 3936 8288
rect 5264 8236 5316 8288
rect 5724 8304 5776 8356
rect 6000 8279 6052 8288
rect 6000 8245 6009 8279
rect 6009 8245 6043 8279
rect 6043 8245 6052 8279
rect 6000 8236 6052 8245
rect 7380 8304 7432 8356
rect 10692 8372 10744 8424
rect 12440 8440 12492 8492
rect 13268 8372 13320 8424
rect 13636 8372 13688 8424
rect 13820 8372 13872 8424
rect 10600 8304 10652 8356
rect 10876 8304 10928 8356
rect 9220 8236 9272 8288
rect 12072 8236 12124 8288
rect 12808 8304 12860 8356
rect 13452 8304 13504 8356
rect 13544 8347 13596 8356
rect 13544 8313 13553 8347
rect 13553 8313 13587 8347
rect 13587 8313 13596 8347
rect 13544 8304 13596 8313
rect 14372 8304 14424 8356
rect 14464 8304 14516 8356
rect 14648 8372 14700 8424
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 14740 8304 14792 8356
rect 14832 8304 14884 8356
rect 15476 8304 15528 8356
rect 15936 8483 15988 8492
rect 15936 8449 15945 8483
rect 15945 8449 15979 8483
rect 15979 8449 15988 8483
rect 15936 8440 15988 8449
rect 15752 8372 15804 8424
rect 16212 8415 16264 8424
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 17224 8372 17276 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 16672 8304 16724 8356
rect 17684 8304 17736 8356
rect 18696 8440 18748 8492
rect 20168 8440 20220 8492
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 18972 8372 19024 8424
rect 19248 8372 19300 8424
rect 21180 8372 21232 8424
rect 22376 8372 22428 8424
rect 24860 8372 24912 8424
rect 20260 8304 20312 8356
rect 13912 8236 13964 8288
rect 18788 8236 18840 8288
rect 18972 8236 19024 8288
rect 19340 8236 19392 8288
rect 20444 8236 20496 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 1860 8032 1912 8084
rect 2412 8032 2464 8084
rect 4988 8032 5040 8084
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 7104 8032 7156 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 1216 7964 1268 8016
rect 1584 7964 1636 8016
rect 3516 7964 3568 8016
rect 3148 7896 3200 7948
rect 9036 8032 9088 8084
rect 9128 8032 9180 8084
rect 10140 8032 10192 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11704 8032 11756 8084
rect 12072 8032 12124 8084
rect 19616 8032 19668 8084
rect 20444 8075 20496 8084
rect 20444 8041 20453 8075
rect 20453 8041 20487 8075
rect 20487 8041 20496 8075
rect 20444 8032 20496 8041
rect 25596 8032 25648 8084
rect 7932 7964 7984 8016
rect 2412 7828 2464 7880
rect 4620 7828 4672 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 9680 7896 9732 7948
rect 1676 7692 1728 7744
rect 4712 7692 4764 7744
rect 8300 7828 8352 7880
rect 9128 7828 9180 7880
rect 9312 7828 9364 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 12256 7964 12308 8016
rect 11244 7896 11296 7948
rect 12440 7896 12492 7948
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 13452 7896 13504 7948
rect 14648 7896 14700 7948
rect 15292 7964 15344 8016
rect 16764 7964 16816 8016
rect 14924 7896 14976 7948
rect 16212 7939 16264 7948
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 16396 7896 16448 7948
rect 19340 7964 19392 8016
rect 24032 7964 24084 8016
rect 10140 7828 10192 7880
rect 8484 7692 8536 7744
rect 8852 7692 8904 7744
rect 12164 7828 12216 7880
rect 13912 7828 13964 7880
rect 19892 7896 19944 7948
rect 20260 7896 20312 7948
rect 22836 7896 22888 7948
rect 24860 7896 24912 7948
rect 17500 7871 17552 7880
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 17592 7828 17644 7880
rect 10968 7692 11020 7744
rect 11796 7692 11848 7744
rect 12532 7692 12584 7744
rect 12808 7735 12860 7744
rect 12808 7701 12817 7735
rect 12817 7701 12851 7735
rect 12851 7701 12860 7735
rect 12808 7692 12860 7701
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 13820 7760 13872 7812
rect 15108 7760 15160 7812
rect 17408 7760 17460 7812
rect 19064 7760 19116 7812
rect 14188 7692 14240 7744
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 16580 7692 16632 7744
rect 19616 7760 19668 7812
rect 19800 7803 19852 7812
rect 19800 7769 19809 7803
rect 19809 7769 19843 7803
rect 19843 7769 19852 7803
rect 19800 7760 19852 7769
rect 19984 7760 20036 7812
rect 22468 7760 22520 7812
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 19340 7692 19392 7744
rect 19708 7692 19760 7744
rect 19892 7735 19944 7744
rect 19892 7701 19901 7735
rect 19901 7701 19935 7735
rect 19935 7701 19944 7735
rect 19892 7692 19944 7701
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 1768 7488 1820 7540
rect 2596 7488 2648 7540
rect 5264 7488 5316 7540
rect 6828 7488 6880 7540
rect 3424 7420 3476 7472
rect 3884 7420 3936 7472
rect 5724 7420 5776 7472
rect 2688 7352 2740 7404
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3976 7352 4028 7404
rect 4068 7352 4120 7404
rect 4344 7352 4396 7404
rect 6000 7352 6052 7404
rect 10324 7488 10376 7540
rect 10416 7488 10468 7540
rect 8576 7420 8628 7472
rect 9496 7420 9548 7472
rect 10968 7488 11020 7540
rect 12624 7488 12676 7540
rect 7472 7352 7524 7404
rect 12072 7352 12124 7404
rect 12348 7352 12400 7404
rect 12440 7352 12492 7404
rect 2320 7216 2372 7268
rect 3148 7284 3200 7336
rect 7012 7284 7064 7336
rect 8760 7284 8812 7336
rect 2872 7216 2924 7268
rect 3516 7216 3568 7268
rect 3976 7259 4028 7268
rect 3976 7225 3985 7259
rect 3985 7225 4019 7259
rect 4019 7225 4028 7259
rect 3976 7216 4028 7225
rect 4988 7216 5040 7268
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 6000 7148 6052 7200
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 10140 7284 10192 7336
rect 11336 7284 11388 7336
rect 10416 7216 10468 7268
rect 12900 7216 12952 7268
rect 9404 7148 9456 7200
rect 11428 7148 11480 7200
rect 11796 7148 11848 7200
rect 11980 7148 12032 7200
rect 12348 7148 12400 7200
rect 15568 7420 15620 7472
rect 16212 7420 16264 7472
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 15936 7352 15988 7404
rect 17408 7420 17460 7472
rect 18236 7420 18288 7472
rect 16764 7352 16816 7404
rect 19248 7352 19300 7404
rect 17408 7284 17460 7336
rect 16028 7216 16080 7268
rect 17132 7216 17184 7268
rect 18604 7284 18656 7336
rect 18880 7284 18932 7336
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 16212 7148 16264 7200
rect 16396 7148 16448 7200
rect 16580 7148 16632 7200
rect 17868 7148 17920 7200
rect 22744 7420 22796 7472
rect 23940 7488 23992 7540
rect 19616 7352 19668 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 22652 7284 22704 7336
rect 24124 7284 24176 7336
rect 23848 7216 23900 7268
rect 25320 7216 25372 7268
rect 19616 7191 19668 7200
rect 19616 7157 19625 7191
rect 19625 7157 19659 7191
rect 19659 7157 19668 7191
rect 19616 7148 19668 7157
rect 22100 7148 22152 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 4620 6944 4672 6996
rect 8944 6987 8996 6996
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 2136 6876 2188 6928
rect 2872 6876 2924 6928
rect 5080 6876 5132 6928
rect 2320 6808 2372 6860
rect 1124 6740 1176 6792
rect 5632 6808 5684 6860
rect 6552 6876 6604 6928
rect 10876 6944 10928 6996
rect 11060 6944 11112 6996
rect 12348 6944 12400 6996
rect 12624 6944 12676 6996
rect 19616 6944 19668 6996
rect 9220 6851 9272 6860
rect 9220 6817 9229 6851
rect 9229 6817 9263 6851
rect 9263 6817 9272 6851
rect 9220 6808 9272 6817
rect 9404 6808 9456 6860
rect 12256 6808 12308 6860
rect 12624 6808 12676 6860
rect 16764 6876 16816 6928
rect 17500 6876 17552 6928
rect 19800 6876 19852 6928
rect 19892 6876 19944 6928
rect 572 6672 624 6724
rect 1308 6672 1360 6724
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6740 4120 6792
rect 4988 6672 5040 6724
rect 5908 6740 5960 6792
rect 6552 6740 6604 6792
rect 6276 6672 6328 6724
rect 8760 6740 8812 6792
rect 8852 6740 8904 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 11980 6740 12032 6792
rect 14004 6808 14056 6860
rect 15752 6808 15804 6860
rect 15936 6808 15988 6860
rect 18512 6808 18564 6860
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 20076 6808 20128 6860
rect 25504 6808 25556 6860
rect 4068 6604 4120 6656
rect 5448 6604 5500 6656
rect 7104 6604 7156 6656
rect 10784 6672 10836 6724
rect 11152 6672 11204 6724
rect 9312 6604 9364 6656
rect 15200 6740 15252 6792
rect 12256 6672 12308 6724
rect 12532 6672 12584 6724
rect 13912 6672 13964 6724
rect 14924 6672 14976 6724
rect 15660 6672 15712 6724
rect 16120 6672 16172 6724
rect 16672 6740 16724 6792
rect 16764 6715 16816 6724
rect 16764 6681 16773 6715
rect 16773 6681 16807 6715
rect 16807 6681 16816 6715
rect 16764 6672 16816 6681
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 12624 6604 12676 6656
rect 13360 6604 13412 6656
rect 14280 6604 14332 6656
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 15016 6604 15068 6613
rect 15292 6604 15344 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 17592 6604 17644 6656
rect 18236 6672 18288 6724
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 18512 6604 18564 6656
rect 20076 6672 20128 6724
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 21916 6715 21968 6724
rect 21916 6681 21925 6715
rect 21925 6681 21959 6715
rect 21959 6681 21968 6715
rect 21916 6672 21968 6681
rect 25044 6672 25096 6724
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 940 6400 992 6452
rect 3148 6400 3200 6452
rect 5172 6332 5224 6384
rect 5264 6332 5316 6384
rect 7656 6332 7708 6384
rect 480 6196 532 6248
rect 2320 6196 2372 6248
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 3884 6196 3936 6248
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 4804 6196 4856 6248
rect 4988 6196 5040 6248
rect 6736 6196 6788 6248
rect 2688 6128 2740 6180
rect 7012 6128 7064 6180
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 8760 6400 8812 6452
rect 11336 6400 11388 6452
rect 11612 6332 11664 6384
rect 11980 6332 12032 6384
rect 13912 6400 13964 6452
rect 14004 6400 14056 6452
rect 14832 6400 14884 6452
rect 15016 6400 15068 6452
rect 17776 6400 17828 6452
rect 12532 6332 12584 6384
rect 14372 6332 14424 6384
rect 15292 6332 15344 6384
rect 15476 6375 15528 6384
rect 15476 6341 15485 6375
rect 15485 6341 15519 6375
rect 15519 6341 15528 6375
rect 15476 6332 15528 6341
rect 16488 6332 16540 6384
rect 9220 6264 9272 6316
rect 9312 6196 9364 6248
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 11244 6196 11296 6248
rect 11796 6196 11848 6248
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 13544 6264 13596 6316
rect 14280 6264 14332 6316
rect 14556 6264 14608 6316
rect 4160 6060 4212 6112
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 6736 6060 6788 6112
rect 6828 6060 6880 6112
rect 8576 6060 8628 6112
rect 8944 6103 8996 6112
rect 8944 6069 8953 6103
rect 8953 6069 8987 6103
rect 8987 6069 8996 6103
rect 8944 6060 8996 6069
rect 9128 6060 9180 6112
rect 11980 6060 12032 6112
rect 12348 6060 12400 6112
rect 13820 6196 13872 6248
rect 15200 6196 15252 6248
rect 15568 6196 15620 6248
rect 15844 6196 15896 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 15936 6128 15988 6180
rect 16396 6264 16448 6316
rect 20444 6400 20496 6452
rect 21732 6400 21784 6452
rect 19248 6332 19300 6384
rect 20260 6264 20312 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 16764 6196 16816 6248
rect 17592 6196 17644 6248
rect 13360 6060 13412 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 17224 6060 17276 6112
rect 17684 6128 17736 6180
rect 18236 6060 18288 6112
rect 19708 6128 19760 6180
rect 21732 6196 21784 6248
rect 19616 6060 19668 6112
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 20536 6060 20588 6112
rect 20628 6060 20680 6112
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 2688 5856 2740 5908
rect 2780 5856 2832 5908
rect 4160 5788 4212 5840
rect 6828 5856 6880 5908
rect 7196 5856 7248 5908
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 11060 5856 11112 5908
rect 11152 5856 11204 5908
rect 12624 5856 12676 5908
rect 13544 5856 13596 5908
rect 13728 5856 13780 5908
rect 4804 5788 4856 5840
rect 7288 5788 7340 5840
rect 7656 5720 7708 5772
rect 7748 5720 7800 5772
rect 2412 5652 2464 5704
rect 2136 5627 2188 5636
rect 2136 5593 2145 5627
rect 2145 5593 2179 5627
rect 2179 5593 2188 5627
rect 2136 5584 2188 5593
rect 3792 5652 3844 5704
rect 5172 5652 5224 5704
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 4160 5584 4212 5636
rect 4620 5584 4672 5636
rect 7564 5652 7616 5704
rect 8944 5652 8996 5704
rect 9588 5584 9640 5636
rect 3608 5516 3660 5568
rect 3792 5516 3844 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 12808 5788 12860 5840
rect 14372 5788 14424 5840
rect 14740 5788 14792 5840
rect 15200 5788 15252 5840
rect 17408 5856 17460 5908
rect 19248 5856 19300 5908
rect 20260 5856 20312 5908
rect 21640 5856 21692 5908
rect 23296 5856 23348 5908
rect 10600 5720 10652 5772
rect 17592 5720 17644 5772
rect 10784 5584 10836 5636
rect 13360 5652 13412 5704
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 18144 5652 18196 5704
rect 18696 5788 18748 5840
rect 19340 5720 19392 5772
rect 20536 5720 20588 5772
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 20812 5652 20864 5704
rect 23572 5720 23624 5772
rect 24032 5720 24084 5772
rect 25320 5720 25372 5772
rect 22836 5652 22888 5704
rect 24492 5652 24544 5704
rect 15108 5584 15160 5636
rect 10968 5559 11020 5568
rect 10968 5525 10977 5559
rect 10977 5525 11011 5559
rect 11011 5525 11020 5559
rect 10968 5516 11020 5525
rect 13360 5516 13412 5568
rect 13912 5516 13964 5568
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 19984 5584 20036 5636
rect 20720 5584 20772 5636
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 20444 5516 20496 5568
rect 22008 5516 22060 5568
rect 24584 5559 24636 5568
rect 24584 5525 24593 5559
rect 24593 5525 24627 5559
rect 24627 5525 24636 5559
rect 24584 5516 24636 5525
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 3976 5312 4028 5364
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 5356 5312 5408 5364
rect 7380 5312 7432 5364
rect 7656 5312 7708 5364
rect 15108 5312 15160 5364
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 16488 5312 16540 5364
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 19616 5312 19668 5364
rect 22100 5312 22152 5364
rect 22744 5312 22796 5364
rect 3608 5176 3660 5228
rect 12164 5244 12216 5296
rect 13360 5287 13412 5296
rect 13360 5253 13369 5287
rect 13369 5253 13403 5287
rect 13403 5253 13412 5287
rect 13360 5244 13412 5253
rect 6092 5176 6144 5228
rect 7104 5176 7156 5228
rect 9312 5176 9364 5228
rect 9956 5176 10008 5228
rect 11612 5219 11664 5228
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 14464 5176 14516 5228
rect 4712 5108 4764 5160
rect 6092 5040 6144 5092
rect 12256 5108 12308 5160
rect 12716 5108 12768 5160
rect 12992 5108 13044 5160
rect 14648 5108 14700 5160
rect 14372 5040 14424 5092
rect 16948 5244 17000 5296
rect 17776 5244 17828 5296
rect 15292 5176 15344 5228
rect 16304 5176 16356 5228
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 18328 5151 18380 5160
rect 18328 5117 18337 5151
rect 18337 5117 18371 5151
rect 18371 5117 18380 5151
rect 18328 5108 18380 5117
rect 14924 5040 14976 5092
rect 21180 5176 21232 5228
rect 4160 4972 4212 5024
rect 4344 4972 4396 5024
rect 8852 4972 8904 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 10324 4972 10376 5024
rect 11612 4972 11664 5024
rect 12808 4972 12860 5024
rect 12992 4972 13044 5024
rect 13452 4972 13504 5024
rect 14832 5015 14884 5024
rect 14832 4981 14841 5015
rect 14841 4981 14875 5015
rect 14875 4981 14884 5015
rect 14832 4972 14884 4981
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 17408 4972 17460 5024
rect 17868 4972 17920 5024
rect 18604 4972 18656 5024
rect 19800 5108 19852 5160
rect 23940 5219 23992 5228
rect 23940 5185 23949 5219
rect 23949 5185 23983 5219
rect 23983 5185 23992 5219
rect 23940 5176 23992 5185
rect 21548 5108 21600 5160
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 7656 4811 7708 4820
rect 7656 4777 7665 4811
rect 7665 4777 7699 4811
rect 7699 4777 7708 4811
rect 7656 4768 7708 4777
rect 8484 4768 8536 4820
rect 9036 4768 9088 4820
rect 9312 4768 9364 4820
rect 15476 4768 15528 4820
rect 15936 4768 15988 4820
rect 17776 4768 17828 4820
rect 19892 4768 19944 4820
rect 9404 4632 9456 4684
rect 14556 4700 14608 4752
rect 14924 4700 14976 4752
rect 16488 4700 16540 4752
rect 19708 4700 19760 4752
rect 1032 4564 1084 4616
rect 1768 4564 1820 4616
rect 2872 4564 2924 4616
rect 3424 4564 3476 4616
rect 8392 4564 8444 4616
rect 8484 4564 8536 4616
rect 9036 4564 9088 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 14832 4632 14884 4684
rect 16028 4632 16080 4684
rect 16120 4632 16172 4684
rect 17868 4632 17920 4684
rect 2872 4471 2924 4480
rect 2872 4437 2881 4471
rect 2881 4437 2915 4471
rect 2915 4437 2924 4471
rect 2872 4428 2924 4437
rect 4068 4428 4120 4480
rect 4436 4428 4488 4480
rect 4804 4428 4856 4480
rect 5356 4539 5408 4548
rect 5356 4505 5365 4539
rect 5365 4505 5399 4539
rect 5399 4505 5408 4539
rect 5356 4496 5408 4505
rect 6644 4428 6696 4480
rect 7656 4428 7708 4480
rect 9220 4496 9272 4548
rect 12808 4564 12860 4616
rect 16488 4564 16540 4616
rect 10324 4428 10376 4480
rect 10508 4428 10560 4480
rect 13728 4428 13780 4480
rect 14648 4428 14700 4480
rect 14740 4428 14792 4480
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20076 4564 20128 4616
rect 18420 4539 18472 4548
rect 18420 4505 18429 4539
rect 18429 4505 18463 4539
rect 18463 4505 18472 4539
rect 18420 4496 18472 4505
rect 19248 4496 19300 4548
rect 20444 4675 20496 4684
rect 20444 4641 20453 4675
rect 20453 4641 20487 4675
rect 20487 4641 20496 4675
rect 20444 4632 20496 4641
rect 20812 4632 20864 4684
rect 21088 4632 21140 4684
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 20812 4496 20864 4548
rect 21180 4496 21232 4548
rect 17316 4428 17368 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 3240 4224 3292 4276
rect 5356 4224 5408 4276
rect 6092 4224 6144 4276
rect 7104 4224 7156 4276
rect 7656 4224 7708 4276
rect 1492 4088 1544 4140
rect 2964 4156 3016 4208
rect 3332 4088 3384 4140
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4988 4088 5040 4140
rect 5632 4088 5684 4140
rect 5908 4088 5960 4140
rect 8760 4156 8812 4208
rect 7012 4088 7064 4140
rect 2412 4020 2464 4072
rect 3516 4063 3568 4072
rect 3516 4029 3525 4063
rect 3525 4029 3559 4063
rect 3559 4029 3568 4063
rect 3516 4020 3568 4029
rect 5264 4020 5316 4072
rect 8944 4088 8996 4140
rect 9772 4224 9824 4276
rect 14372 4224 14424 4276
rect 14464 4224 14516 4276
rect 9680 4156 9732 4208
rect 14280 4156 14332 4208
rect 15844 4224 15896 4276
rect 16028 4224 16080 4276
rect 17132 4224 17184 4276
rect 15660 4156 15712 4208
rect 18788 4224 18840 4276
rect 19248 4224 19300 4276
rect 24308 4224 24360 4276
rect 10140 4088 10192 4140
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 10968 4088 11020 4140
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 13452 4088 13504 4140
rect 10048 4020 10100 4072
rect 2964 3952 3016 4004
rect 11888 4020 11940 4072
rect 14648 4020 14700 4072
rect 16396 4131 16448 4140
rect 16396 4097 16405 4131
rect 16405 4097 16439 4131
rect 16439 4097 16448 4131
rect 16396 4088 16448 4097
rect 18512 4156 18564 4208
rect 19892 4156 19944 4208
rect 21364 4156 21416 4208
rect 19616 4088 19668 4140
rect 20260 4088 20312 4140
rect 21548 4088 21600 4140
rect 22192 4131 22244 4140
rect 22192 4097 22201 4131
rect 22201 4097 22235 4131
rect 22235 4097 22244 4131
rect 22192 4088 22244 4097
rect 22836 4088 22888 4140
rect 23572 4088 23624 4140
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 23940 4088 23992 4140
rect 24952 4088 25004 4140
rect 17592 4063 17644 4072
rect 3792 3884 3844 3936
rect 4436 3884 4488 3936
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6460 3884 6512 3936
rect 7748 3884 7800 3936
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 9680 3884 9732 3936
rect 10140 3884 10192 3936
rect 12624 3884 12676 3936
rect 12716 3884 12768 3936
rect 17592 4029 17601 4063
rect 17601 4029 17635 4063
rect 17635 4029 17644 4063
rect 17592 4020 17644 4029
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 16028 3927 16080 3936
rect 16028 3893 16037 3927
rect 16037 3893 16071 3927
rect 16071 3893 16080 3927
rect 16028 3884 16080 3893
rect 16764 3884 16816 3936
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 19708 4020 19760 4072
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 20720 4020 20772 4072
rect 20812 4020 20864 4072
rect 21456 4020 21508 4072
rect 21364 3952 21416 4004
rect 19708 3884 19760 3936
rect 19984 3927 20036 3936
rect 19984 3893 19993 3927
rect 19993 3893 20027 3927
rect 20027 3893 20036 3927
rect 19984 3884 20036 3893
rect 20168 3884 20220 3936
rect 20352 3884 20404 3936
rect 21640 3884 21692 3936
rect 24952 3884 25004 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 2504 3612 2556 3664
rect 3424 3680 3476 3732
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 4528 3680 4580 3732
rect 7012 3680 7064 3732
rect 7380 3680 7432 3732
rect 5724 3612 5776 3664
rect 6000 3612 6052 3664
rect 7104 3612 7156 3664
rect 664 3476 716 3528
rect 1400 3476 1452 3528
rect 1860 3476 1912 3528
rect 2044 3476 2096 3528
rect 3240 3544 3292 3596
rect 3792 3544 3844 3596
rect 4344 3544 4396 3596
rect 10692 3680 10744 3732
rect 11980 3680 12032 3732
rect 12624 3680 12676 3732
rect 15936 3680 15988 3732
rect 17316 3680 17368 3732
rect 18328 3680 18380 3732
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3424 3476 3476 3528
rect 4160 3476 4212 3528
rect 2964 3408 3016 3460
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 16764 3612 16816 3664
rect 16948 3612 17000 3664
rect 18420 3612 18472 3664
rect 12716 3544 12768 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 1400 3340 1452 3392
rect 11704 3408 11756 3460
rect 12072 3408 12124 3460
rect 13452 3476 13504 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 15752 3476 15804 3528
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 18696 3476 18748 3528
rect 15108 3408 15160 3460
rect 23848 3680 23900 3732
rect 24216 3723 24268 3732
rect 24216 3689 24225 3723
rect 24225 3689 24259 3723
rect 24259 3689 24268 3723
rect 24216 3680 24268 3689
rect 23296 3655 23348 3664
rect 23296 3621 23305 3655
rect 23305 3621 23339 3655
rect 23339 3621 23348 3655
rect 23296 3612 23348 3621
rect 23664 3655 23716 3664
rect 23664 3621 23673 3655
rect 23673 3621 23707 3655
rect 23707 3621 23716 3655
rect 23664 3612 23716 3621
rect 19708 3544 19760 3596
rect 20444 3544 20496 3596
rect 20720 3544 20772 3596
rect 22560 3544 22612 3596
rect 21180 3476 21232 3528
rect 21640 3519 21692 3528
rect 21640 3485 21649 3519
rect 21649 3485 21683 3519
rect 21683 3485 21692 3519
rect 21640 3476 21692 3485
rect 23296 3476 23348 3528
rect 24308 3476 24360 3528
rect 24492 3476 24544 3528
rect 19708 3451 19760 3460
rect 19708 3417 19717 3451
rect 19717 3417 19751 3451
rect 19751 3417 19760 3451
rect 19708 3408 19760 3417
rect 22008 3408 22060 3460
rect 24216 3408 24268 3460
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8300 3340 8352 3392
rect 9404 3340 9456 3392
rect 11796 3340 11848 3392
rect 17132 3340 17184 3392
rect 17592 3340 17644 3392
rect 23480 3340 23532 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 1216 3136 1268 3188
rect 1676 3111 1728 3120
rect 1676 3077 1685 3111
rect 1685 3077 1719 3111
rect 1719 3077 1728 3111
rect 1676 3068 1728 3077
rect 1860 3111 1912 3120
rect 1860 3077 1869 3111
rect 1869 3077 1903 3111
rect 1903 3077 1912 3111
rect 1860 3068 1912 3077
rect 3240 3136 3292 3188
rect 3792 3136 3844 3188
rect 3884 3136 3936 3188
rect 4620 3136 4672 3188
rect 5724 3136 5776 3188
rect 6276 3136 6328 3188
rect 6644 3136 6696 3188
rect 6828 3136 6880 3188
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 13360 3136 13412 3188
rect 18788 3136 18840 3188
rect 20720 3136 20772 3188
rect 7380 3068 7432 3120
rect 7656 3068 7708 3120
rect 8760 3068 8812 3120
rect 9956 3068 10008 3120
rect 23388 3068 23440 3120
rect 2688 3000 2740 3052
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 6092 3000 6144 3052
rect 2872 2932 2924 2984
rect 756 2796 808 2848
rect 6184 2932 6236 2984
rect 6920 3000 6972 3052
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 8576 2932 8628 2984
rect 9956 2932 10008 2984
rect 11428 2932 11480 2984
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 10692 2864 10744 2916
rect 11520 2864 11572 2916
rect 12072 2932 12124 2984
rect 12532 2932 12584 2984
rect 13360 3000 13412 3052
rect 16580 3000 16632 3052
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 21272 3000 21324 3052
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 23848 3043 23900 3052
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 16120 2864 16172 2916
rect 16212 2864 16264 2916
rect 19524 2932 19576 2984
rect 21456 2932 21508 2984
rect 3792 2796 3844 2848
rect 8300 2796 8352 2848
rect 18236 2796 18288 2848
rect 19892 2796 19944 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 1492 2635 1544 2644
rect 1492 2601 1501 2635
rect 1501 2601 1535 2635
rect 1535 2601 1544 2635
rect 1492 2592 1544 2601
rect 3424 2592 3476 2644
rect 3516 2592 3568 2644
rect 13360 2592 13412 2644
rect 2688 2524 2740 2576
rect 3700 2456 3752 2508
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 3332 2388 3384 2440
rect 3608 2388 3660 2440
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 5724 2456 5776 2508
rect 8484 2456 8536 2508
rect 9036 2456 9088 2508
rect 12440 2456 12492 2508
rect 14372 2456 14424 2508
rect 15108 2456 15160 2508
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5816 2388 5868 2440
rect 5908 2388 5960 2440
rect 7288 2320 7340 2372
rect 848 2252 900 2304
rect 7748 2252 7800 2304
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 10968 2363 11020 2372
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 15568 2320 15620 2372
rect 15936 2320 15988 2372
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 14924 2252 14976 2304
rect 16028 2252 16080 2304
rect 17132 2388 17184 2440
rect 17684 2592 17736 2644
rect 19064 2592 19116 2644
rect 22284 2592 22336 2644
rect 22376 2592 22428 2644
rect 23204 2592 23256 2644
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 24492 2592 24544 2644
rect 24584 2592 24636 2644
rect 18972 2456 19024 2508
rect 24216 2567 24268 2576
rect 24216 2533 24225 2567
rect 24225 2533 24259 2567
rect 24259 2533 24268 2567
rect 24216 2524 24268 2533
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 16672 2320 16724 2372
rect 21824 2388 21876 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 21088 2295 21140 2304
rect 21088 2261 21097 2295
rect 21097 2261 21131 2295
rect 21131 2261 21140 2295
rect 21088 2252 21140 2261
rect 21272 2295 21324 2304
rect 21272 2261 21281 2295
rect 21281 2261 21315 2295
rect 21315 2261 21324 2295
rect 21272 2252 21324 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 7564 2048 7616 2100
rect 8116 2048 8168 2100
rect 3424 1980 3476 2032
rect 11796 1980 11848 2032
rect 7196 1912 7248 1964
rect 19800 1912 19852 1964
rect 2412 1844 2464 1896
rect 14096 1844 14148 1896
rect 4620 1776 4672 1828
rect 10324 1776 10376 1828
rect 10968 1776 11020 1828
rect 22192 1776 22244 1828
rect 5356 1708 5408 1760
rect 13912 1708 13964 1760
rect 2136 1640 2188 1692
rect 17500 1640 17552 1692
rect 5264 1572 5316 1624
rect 9772 1572 9824 1624
rect 9496 1504 9548 1556
rect 24584 1504 24636 1556
rect 9312 1436 9364 1488
rect 17224 1436 17276 1488
rect 1768 1368 1820 1420
rect 9588 1368 9640 1420
rect 7932 1300 7984 1352
rect 24400 1300 24452 1352
rect 8668 1232 8720 1284
rect 21272 1232 21324 1284
rect 6460 1164 6512 1216
rect 20076 1164 20128 1216
rect 4160 1096 4212 1148
rect 18880 1096 18932 1148
rect 8300 1028 8352 1080
rect 21088 1028 21140 1080
rect 7840 960 7892 1012
rect 19616 960 19668 1012
rect 7656 892 7708 944
rect 20904 892 20956 944
rect 7472 824 7524 876
rect 19708 824 19760 876
rect 4344 144 4396 196
rect 12440 144 12492 196
rect 6184 76 6236 128
rect 24216 76 24268 128
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 3896 56222 4108 56250
rect 1044 53650 1072 56200
rect 2424 54126 2452 56200
rect 3804 56114 3832 56200
rect 3896 56114 3924 56222
rect 3804 56086 3924 56114
rect 3884 54188 3936 54194
rect 3884 54130 3936 54136
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3896 53242 3924 54130
rect 4080 54126 4108 56222
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 6656 56222 6868 56250
rect 4068 54120 4120 54126
rect 4068 54062 4120 54068
rect 5184 53650 5212 56200
rect 6564 56114 6592 56200
rect 6656 56114 6684 56222
rect 6564 56086 6684 56114
rect 6840 54210 6868 56222
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 10796 56222 11008 56250
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 6552 54188 6604 54194
rect 6552 54130 6604 54136
rect 6736 54188 6788 54194
rect 6840 54182 6960 54210
rect 6736 54130 6788 54136
rect 5172 53644 5224 53650
rect 5172 53586 5224 53592
rect 5540 53508 5592 53514
rect 5540 53450 5592 53456
rect 3884 53236 3936 53242
rect 3884 53178 3936 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 5552 50726 5580 53450
rect 6564 53242 6592 54130
rect 6552 53236 6604 53242
rect 6552 53178 6604 53184
rect 6748 52154 6776 54130
rect 6932 54126 6960 54182
rect 6920 54120 6972 54126
rect 6920 54062 6972 54068
rect 7656 53576 7708 53582
rect 7656 53518 7708 53524
rect 7668 52698 7696 53518
rect 7748 53032 7800 53038
rect 7748 52974 7800 52980
rect 7656 52692 7708 52698
rect 7656 52634 7708 52640
rect 6736 52148 6788 52154
rect 6736 52090 6788 52096
rect 7760 51066 7788 52974
rect 7852 52630 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 8852 53100 8904 53106
rect 8852 53042 8904 53048
rect 7840 52624 7892 52630
rect 7840 52566 7892 52572
rect 8392 52624 8444 52630
rect 8392 52566 8444 52572
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7748 51060 7800 51066
rect 7748 51002 7800 51008
rect 5540 50720 5592 50726
rect 5540 50662 5592 50668
rect 6828 50720 6880 50726
rect 6828 50662 6880 50668
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 6840 50386 6868 50662
rect 6828 50380 6880 50386
rect 6828 50322 6880 50328
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 7760 48822 7788 51002
rect 8300 50380 8352 50386
rect 8300 50322 8352 50328
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7748 48816 7800 48822
rect 7748 48758 7800 48764
rect 8208 48816 8260 48822
rect 8208 48758 8260 48764
rect 7748 48680 7800 48686
rect 7748 48622 7800 48628
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 7760 39098 7788 48622
rect 8220 48142 8248 48758
rect 8312 48278 8340 50322
rect 8404 48686 8432 52566
rect 8864 48890 8892 53042
rect 8852 48884 8904 48890
rect 8852 48826 8904 48832
rect 8392 48680 8444 48686
rect 8392 48622 8444 48628
rect 8300 48272 8352 48278
rect 8300 48214 8352 48220
rect 8576 48204 8628 48210
rect 8576 48146 8628 48152
rect 8208 48136 8260 48142
rect 8208 48078 8260 48084
rect 7840 48068 7892 48074
rect 7840 48010 7892 48016
rect 7852 47462 7880 48010
rect 8588 48006 8616 48146
rect 8576 48000 8628 48006
rect 8576 47942 8628 47948
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7840 47456 7892 47462
rect 7840 47398 7892 47404
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 8588 44946 8616 47942
rect 8864 47734 8892 48826
rect 9128 48136 9180 48142
rect 9128 48078 9180 48084
rect 8852 47728 8904 47734
rect 8852 47670 8904 47676
rect 8760 47524 8812 47530
rect 8760 47466 8812 47472
rect 8576 44940 8628 44946
rect 8576 44882 8628 44888
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7748 39092 7800 39098
rect 7748 39034 7800 39040
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 8772 35834 8800 47466
rect 9140 47258 9168 48078
rect 9324 47598 9352 56200
rect 10704 56114 10732 56200
rect 10796 56114 10824 56222
rect 10704 56086 10824 56114
rect 9588 52488 9640 52494
rect 9588 52430 9640 52436
rect 9600 47598 9628 52430
rect 10784 52012 10836 52018
rect 10784 51954 10836 51960
rect 10140 48544 10192 48550
rect 10140 48486 10192 48492
rect 9312 47592 9364 47598
rect 9312 47534 9364 47540
rect 9588 47592 9640 47598
rect 9588 47534 9640 47540
rect 9128 47252 9180 47258
rect 9128 47194 9180 47200
rect 9600 47190 9628 47534
rect 9588 47184 9640 47190
rect 9588 47126 9640 47132
rect 9312 45960 9364 45966
rect 9312 45902 9364 45908
rect 9036 45416 9088 45422
rect 9036 45358 9088 45364
rect 8852 38956 8904 38962
rect 8852 38898 8904 38904
rect 8760 35828 8812 35834
rect 8760 35770 8812 35776
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 4342 29064 4398 29073
rect 4342 28999 4398 29008
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 4252 26920 4304 26926
rect 4252 26862 4304 26868
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3712 19310 3740 21830
rect 3974 19952 4030 19961
rect 3974 19887 4030 19896
rect 3988 19378 4016 19887
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 4264 19310 4292 26862
rect 4356 19922 4384 28999
rect 5538 27432 5594 27441
rect 5538 27367 5594 27376
rect 5552 23474 5580 27367
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6840 26382 6868 26726
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 7484 24818 7512 25638
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6472 23866 6500 24142
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6932 23730 6960 24006
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 7196 23656 7248 23662
rect 7194 23624 7196 23633
rect 7248 23624 7250 23633
rect 7194 23559 7250 23568
rect 5460 23446 5580 23474
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 4356 19514 4384 19858
rect 4620 19848 4672 19854
rect 4618 19816 4620 19825
rect 4672 19816 4674 19825
rect 4618 19751 4674 19760
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 1306 17776 1362 17785
rect 1306 17711 1362 17720
rect 664 16108 716 16114
rect 664 16050 716 16056
rect 572 15700 624 15706
rect 572 15642 624 15648
rect 480 15360 532 15366
rect 480 15302 532 15308
rect 492 6254 520 15302
rect 584 6730 612 15642
rect 572 6724 624 6730
rect 572 6666 624 6672
rect 480 6248 532 6254
rect 480 6190 532 6196
rect 676 3534 704 16050
rect 848 16040 900 16046
rect 848 15982 900 15988
rect 756 15496 808 15502
rect 756 15438 808 15444
rect 664 3528 716 3534
rect 664 3470 716 3476
rect 768 2854 796 15438
rect 756 2848 808 2854
rect 756 2790 808 2796
rect 860 2310 888 15982
rect 1032 15428 1084 15434
rect 1032 15370 1084 15376
rect 940 14884 992 14890
rect 940 14826 992 14832
rect 952 6458 980 14826
rect 940 6452 992 6458
rect 940 6394 992 6400
rect 1044 4622 1072 15370
rect 1216 14952 1268 14958
rect 1216 14894 1268 14900
rect 1124 12640 1176 12646
rect 1124 12582 1176 12588
rect 1136 8294 1164 12582
rect 1124 8288 1176 8294
rect 1124 8230 1176 8236
rect 1228 8106 1256 14894
rect 1320 9450 1348 17711
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1766 15600 1822 15609
rect 1766 15535 1822 15544
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 10742 1440 14214
rect 1400 10736 1452 10742
rect 1400 10678 1452 10684
rect 1412 10130 1440 10678
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1400 9988 1452 9994
rect 1400 9930 1452 9936
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1136 8078 1256 8106
rect 1136 6798 1164 8078
rect 1216 8016 1268 8022
rect 1216 7958 1268 7964
rect 1124 6792 1176 6798
rect 1124 6734 1176 6740
rect 1032 4616 1084 4622
rect 1032 4558 1084 4564
rect 1228 3194 1256 7958
rect 1412 6914 1440 9930
rect 1504 9586 1532 14758
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1596 8906 1624 13126
rect 1688 8974 1716 14758
rect 1780 14074 1808 15535
rect 2056 15366 2084 16186
rect 2504 15972 2556 15978
rect 2504 15914 2556 15920
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2044 15360 2096 15366
rect 2042 15328 2044 15337
rect 2096 15328 2098 15337
rect 2042 15263 2098 15272
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1872 13977 1900 14214
rect 1858 13968 1914 13977
rect 1858 13903 1914 13912
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1780 12753 1808 13262
rect 1766 12744 1822 12753
rect 1766 12679 1768 12688
rect 1820 12679 1822 12688
rect 1768 12650 1820 12656
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 7721 1532 8774
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8022 1624 8434
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1676 7744 1728 7750
rect 1490 7712 1546 7721
rect 1676 7686 1728 7692
rect 1490 7647 1546 7656
rect 1412 6886 1624 6914
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 5545 1348 6666
rect 1306 5536 1362 5545
rect 1306 5471 1362 5480
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1412 3398 1440 3470
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1216 3188 1268 3194
rect 1216 3130 1268 3136
rect 1412 2530 1440 3334
rect 1504 2650 1532 4082
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1412 2502 1532 2530
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 1504 800 1532 2502
rect 1490 0 1546 800
rect 1596 762 1624 6886
rect 1688 4593 1716 7686
rect 1780 7546 1808 11086
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 10810 1900 10950
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1860 9512 1912 9518
rect 1858 9480 1860 9489
rect 1912 9480 1914 9489
rect 1858 9415 1914 9424
rect 1964 8498 1992 14758
rect 2056 14414 2084 14758
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 14249 2084 14350
rect 2042 14240 2098 14249
rect 2042 14175 2098 14184
rect 2148 13870 2176 15846
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 12345 2176 13806
rect 2134 12336 2190 12345
rect 2134 12271 2190 12280
rect 2136 12232 2188 12238
rect 2134 12200 2136 12209
rect 2188 12200 2190 12209
rect 2134 12135 2190 12144
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 10985 2084 11698
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2042 10976 2098 10985
rect 2042 10911 2098 10920
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2056 9761 2084 10542
rect 2042 9752 2098 9761
rect 2042 9687 2098 9696
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1950 8392 2006 8401
rect 1950 8327 2006 8336
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1768 4616 1820 4622
rect 1674 4584 1730 4593
rect 1768 4558 1820 4564
rect 1674 4519 1730 4528
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1688 3126 1716 3975
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1780 1426 1808 4558
rect 1872 3534 1900 8026
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1858 3224 1914 3233
rect 1858 3159 1914 3168
rect 1872 3126 1900 3159
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1964 2446 1992 8327
rect 2056 3534 2084 8910
rect 2148 6934 2176 11494
rect 2240 9674 2268 15302
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 2332 13326 2360 14486
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2240 9646 2360 9674
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2148 1698 2176 5578
rect 2136 1692 2188 1698
rect 2136 1634 2188 1640
rect 1768 1420 1820 1426
rect 1768 1362 1820 1368
rect 1780 870 1900 898
rect 1780 762 1808 870
rect 1872 800 1900 870
rect 2240 800 2268 9522
rect 2332 9450 2360 9646
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2332 7698 2360 9386
rect 2424 9042 2452 15302
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 8090 2452 8978
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2410 7984 2466 7993
rect 2410 7919 2466 7928
rect 2424 7886 2452 7919
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2332 7670 2452 7698
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 6866 2360 7210
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2332 1737 2360 6190
rect 2424 5710 2452 7670
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2424 1902 2452 4014
rect 2516 3670 2544 15914
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 13841 2636 14758
rect 2700 14414 2728 16934
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2792 13938 2820 19110
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 4264 18766 4292 19246
rect 4252 18760 4304 18766
rect 4066 18728 4122 18737
rect 4252 18702 4304 18708
rect 4066 18663 4122 18672
rect 4080 18630 4108 18663
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4540 18358 4568 18566
rect 4528 18352 4580 18358
rect 4724 18306 4752 21490
rect 5170 21448 5226 21457
rect 5170 21383 5226 21392
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 20398 5120 20742
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5092 19417 5120 20334
rect 5078 19408 5134 19417
rect 5078 19343 5134 19352
rect 4528 18294 4580 18300
rect 4632 18278 4752 18306
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 3422 15736 3478 15745
rect 3422 15671 3478 15680
rect 3436 15638 3464 15671
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2594 13832 2650 13841
rect 2594 13767 2650 13776
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2608 10826 2636 13466
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2700 11082 2728 11698
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2792 11014 2820 11086
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2608 10798 2820 10826
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2700 10169 2728 10406
rect 2686 10160 2742 10169
rect 2686 10095 2742 10104
rect 2686 9888 2742 9897
rect 2686 9823 2742 9832
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 7546 2636 9318
rect 2700 8974 2728 9823
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2792 8566 2820 10798
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2686 8392 2742 8401
rect 2686 8327 2688 8336
rect 2740 8327 2742 8336
rect 2688 8298 2740 8304
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2700 6304 2728 7346
rect 2608 6276 2728 6304
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2608 3618 2636 6276
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 5914 2728 6122
rect 2792 5914 2820 7346
rect 2884 7274 2912 15302
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3252 14929 3280 14962
rect 3238 14920 3294 14929
rect 3238 14855 3294 14864
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3238 11112 3294 11121
rect 3238 11047 3240 11056
rect 3292 11047 3294 11056
rect 3240 11018 3292 11024
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 3238 10024 3294 10033
rect 3238 9959 3240 9968
rect 3292 9959 3294 9968
rect 3240 9930 3292 9936
rect 3240 9648 3292 9654
rect 3238 9616 3240 9625
rect 3292 9616 3294 9625
rect 3238 9551 3294 9560
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8634 3188 8774
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3160 7342 3188 7890
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2884 4622 2912 6870
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3160 6254 3188 6394
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4185 2912 4422
rect 3252 4282 3280 4655
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 2964 4208 3016 4214
rect 2870 4176 2926 4185
rect 2964 4150 3016 4156
rect 2870 4111 2926 4120
rect 2870 4040 2926 4049
rect 2976 4010 3004 4150
rect 3344 4146 3372 15506
rect 3436 14906 3464 15574
rect 3436 14878 3556 14906
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 13705 3464 14758
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 10062 3464 13194
rect 3528 11626 3556 14878
rect 3620 12986 3648 16934
rect 3804 16182 3832 18022
rect 4526 17912 4582 17921
rect 4526 17847 4582 17856
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 4066 16008 4122 16017
rect 4066 15943 4122 15952
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3606 12472 3662 12481
rect 3606 12407 3662 12416
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3620 10690 3648 12407
rect 3528 10662 3648 10690
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3528 9110 3556 10662
rect 3608 10600 3660 10606
rect 3606 10568 3608 10577
rect 3660 10568 3662 10577
rect 3606 10503 3662 10512
rect 3606 10432 3662 10441
rect 3606 10367 3662 10376
rect 3516 9104 3568 9110
rect 3422 9072 3478 9081
rect 3516 9046 3568 9052
rect 3422 9007 3478 9016
rect 3436 8974 3464 9007
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 7478 3464 8910
rect 3514 8120 3570 8129
rect 3514 8055 3570 8064
rect 3528 8022 3556 8055
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 4622 3464 7142
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3528 4162 3556 7210
rect 3620 5574 3648 10367
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3436 4134 3556 4162
rect 2870 3975 2926 3984
rect 2964 4004 3016 4010
rect 2516 3482 2544 3606
rect 2608 3590 2728 3618
rect 2700 3482 2728 3590
rect 2884 3534 2912 3975
rect 2964 3946 3016 3952
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 2872 3528 2924 3534
rect 2516 3454 2636 3482
rect 2700 3454 2820 3482
rect 2872 3470 2924 3476
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2318 1728 2374 1737
rect 2318 1663 2374 1672
rect 2608 800 2636 3454
rect 2686 3360 2742 3369
rect 2686 3295 2742 3304
rect 2700 3058 2728 3295
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2792 2938 2820 3454
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2700 2910 2820 2938
rect 2872 2984 2924 2990
rect 2976 2972 3004 3402
rect 3252 3194 3280 3538
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2924 2944 3004 2972
rect 2872 2926 2924 2932
rect 2700 2582 2728 2910
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2884 2530 2912 2926
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2530 3372 4082
rect 3436 3738 3464 4134
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3436 2650 3464 3470
rect 3528 2650 3556 4014
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 2884 2502 3004 2530
rect 3344 2502 3464 2530
rect 2976 800 3004 2502
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3344 800 3372 2382
rect 3436 2038 3464 2502
rect 3620 2446 3648 5170
rect 3712 2514 3740 15302
rect 3896 15026 3924 15302
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3790 14784 3846 14793
rect 3790 14719 3846 14728
rect 3804 13977 3832 14719
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3896 14414 3924 14554
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3896 13190 3924 13874
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12646 3832 12786
rect 3792 12640 3844 12646
rect 3790 12608 3792 12617
rect 3844 12608 3846 12617
rect 3790 12543 3846 12552
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 8566 3832 12038
rect 3896 11762 3924 12922
rect 3988 12186 4016 15370
rect 4080 14618 4108 15943
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4080 13977 4108 14282
rect 4066 13968 4122 13977
rect 4066 13903 4122 13912
rect 4172 13326 4200 15846
rect 4250 15464 4306 15473
rect 4250 15399 4252 15408
rect 4304 15399 4306 15408
rect 4252 15370 4304 15376
rect 4356 14958 4384 16594
rect 4448 16250 4476 17070
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4448 15881 4476 16186
rect 4434 15872 4490 15881
rect 4434 15807 4490 15816
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4448 15162 4476 15438
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4540 14804 4568 17847
rect 4356 14776 4568 14804
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4264 13433 4292 13874
rect 4250 13424 4306 13433
rect 4250 13359 4306 13368
rect 4264 13326 4292 13359
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4066 12336 4122 12345
rect 4066 12271 4068 12280
rect 4120 12271 4122 12280
rect 4068 12242 4120 12248
rect 4252 12232 4304 12238
rect 3988 12158 4108 12186
rect 4252 12174 4304 12180
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11801 4016 12038
rect 3974 11792 4030 11801
rect 3884 11756 3936 11762
rect 3974 11727 3976 11736
rect 3884 11698 3936 11704
rect 4028 11727 4030 11736
rect 3976 11698 4028 11704
rect 4080 11642 4108 12158
rect 3988 11614 4108 11642
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3896 8378 3924 11290
rect 3988 8945 4016 11614
rect 4264 11558 4292 12174
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 9382 4108 11086
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3974 8936 4030 8945
rect 3974 8871 4030 8880
rect 3976 8832 4028 8838
rect 4080 8809 4108 9046
rect 3976 8774 4028 8780
rect 4066 8800 4122 8809
rect 3804 8350 3924 8378
rect 3804 5710 3832 8350
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7478 3924 8230
rect 3988 8129 4016 8774
rect 4066 8735 4122 8744
rect 4172 8566 4200 11494
rect 4356 11150 4384 14776
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4448 10996 4476 14486
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12442 4568 13262
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4356 10968 4476 10996
rect 4250 10296 4306 10305
rect 4250 10231 4306 10240
rect 4264 10198 4292 10231
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 4080 7410 4108 8434
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3988 7274 4016 7346
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3976 6792 4028 6798
rect 4068 6792 4120 6798
rect 3976 6734 4028 6740
rect 4066 6760 4068 6769
rect 4120 6760 4122 6769
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 3942 3832 5510
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3804 3602 3832 3674
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3896 3194 3924 6190
rect 3988 5370 4016 6734
rect 4066 6695 4122 6704
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4080 4706 4108 6598
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5846 4200 6054
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4158 5672 4214 5681
rect 4158 5607 4160 5616
rect 4212 5607 4214 5616
rect 4160 5578 4212 5584
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3988 4678 4108 4706
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3804 2938 3832 3130
rect 3882 3088 3938 3097
rect 3882 3023 3884 3032
rect 3936 3023 3938 3032
rect 3884 2994 3936 3000
rect 3804 2910 3924 2938
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 3804 1442 3832 2790
rect 3712 1414 3832 1442
rect 3896 1442 3924 2910
rect 3988 2446 4016 4678
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4080 4321 4108 4422
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4172 3534 4200 4966
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4264 2774 4292 9522
rect 4356 7528 4384 10968
rect 4540 9654 4568 11562
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4448 7993 4476 9590
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4434 7984 4490 7993
rect 4434 7919 4490 7928
rect 4356 7500 4476 7528
rect 4342 7440 4398 7449
rect 4342 7375 4344 7384
rect 4396 7375 4398 7384
rect 4344 7346 4396 7352
rect 4344 6248 4396 6254
rect 4342 6216 4344 6225
rect 4396 6216 4398 6225
rect 4342 6151 4398 6160
rect 4356 5030 4384 6151
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4448 4486 4476 7500
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4172 2746 4292 2774
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 3896 1414 4108 1442
rect 3712 800 3740 1414
rect 4080 800 4108 1414
rect 4172 1154 4200 2746
rect 4160 1148 4212 1154
rect 4160 1090 4212 1096
rect 1596 734 1808 762
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4356 202 4384 3538
rect 4448 800 4476 3878
rect 4540 3738 4568 9318
rect 4632 8974 4660 18278
rect 4712 18216 4764 18222
rect 4710 18184 4712 18193
rect 4764 18184 4766 18193
rect 4710 18119 4766 18128
rect 4894 17232 4950 17241
rect 4894 17167 4950 17176
rect 4710 17096 4766 17105
rect 4710 17031 4766 17040
rect 4724 12374 4752 17031
rect 4908 16114 4936 17167
rect 4986 16144 5042 16153
rect 4896 16108 4948 16114
rect 4986 16079 5042 16088
rect 4896 16050 4948 16056
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11286 4752 12038
rect 4816 11898 4844 12922
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10742 4752 10950
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4724 7886 4752 9114
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4632 7002 4660 7822
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4632 3777 4660 5578
rect 4724 5166 4752 7686
rect 4816 6254 4844 11018
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 8650 4936 10950
rect 5000 10538 5028 16079
rect 5078 15464 5134 15473
rect 5078 15399 5134 15408
rect 5092 13138 5120 15399
rect 5184 14550 5212 21383
rect 5354 20088 5410 20097
rect 5354 20023 5410 20032
rect 5368 17338 5396 20023
rect 5460 17746 5488 23446
rect 6274 23216 6330 23225
rect 6274 23151 6330 23160
rect 6288 23118 6316 23151
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 6276 22228 6328 22234
rect 6276 22170 6328 22176
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6012 19514 6040 20402
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6182 19272 6238 19281
rect 6000 19236 6052 19242
rect 6182 19207 6238 19216
rect 6000 19178 6052 19184
rect 6012 18902 6040 19178
rect 6000 18896 6052 18902
rect 5722 18864 5778 18873
rect 6000 18838 6052 18844
rect 5722 18799 5778 18808
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5368 15706 5396 17138
rect 5644 16794 5672 17614
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5552 16250 5580 16662
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5460 14958 5488 15098
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 5262 14376 5318 14385
rect 5262 14311 5264 14320
rect 5316 14311 5318 14320
rect 5264 14282 5316 14288
rect 5736 14090 5764 18799
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 18426 6040 18702
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6090 17640 6146 17649
rect 6090 17575 6146 17584
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5644 14062 5764 14090
rect 5644 13462 5672 14062
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5170 13288 5226 13297
rect 5170 13223 5172 13232
rect 5224 13223 5226 13232
rect 5448 13252 5500 13258
rect 5172 13194 5224 13200
rect 5448 13194 5500 13200
rect 5356 13184 5408 13190
rect 5092 13110 5212 13138
rect 5356 13126 5408 13132
rect 5078 12880 5134 12889
rect 5078 12815 5080 12824
rect 5132 12815 5134 12824
rect 5080 12786 5132 12792
rect 5092 11898 5120 12786
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 9920 5040 9926
rect 4986 9888 4988 9897
rect 5040 9888 5042 9897
rect 4986 9823 5042 9832
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8809 5028 9318
rect 4986 8800 5042 8809
rect 4986 8735 5042 8744
rect 4908 8622 5028 8650
rect 5000 8378 5028 8622
rect 4908 8350 5028 8378
rect 4908 7970 4936 8350
rect 4986 8256 5042 8265
rect 4986 8191 5042 8200
rect 5000 8090 5028 8191
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4908 7942 5028 7970
rect 4894 7712 4950 7721
rect 4894 7647 4950 7656
rect 4908 7206 4936 7647
rect 5000 7274 5028 7942
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 7200 4948 7206
rect 4894 7168 4896 7177
rect 4948 7168 4950 7177
rect 4894 7103 4950 7112
rect 4894 7032 4950 7041
rect 4894 6967 4950 6976
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5846 4844 6054
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4146 4844 4422
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4618 3768 4674 3777
rect 4528 3732 4580 3738
rect 4618 3703 4674 3712
rect 4528 3674 4580 3680
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4632 1834 4660 3130
rect 4908 3058 4936 6967
rect 5092 6934 5120 10406
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4988 6724 5040 6730
rect 5040 6684 5120 6712
rect 4988 6666 5040 6672
rect 5092 6361 5120 6684
rect 5184 6390 5212 13110
rect 5368 12850 5396 13126
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5460 12714 5488 13194
rect 5552 12753 5580 13330
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5538 12744 5594 12753
rect 5448 12708 5500 12714
rect 5644 12714 5672 13262
rect 5538 12679 5594 12688
rect 5632 12708 5684 12714
rect 5448 12650 5500 12656
rect 5632 12650 5684 12656
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5630 12608 5686 12617
rect 5368 11762 5396 12582
rect 5630 12543 5686 12552
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5276 9722 5304 10746
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5264 8968 5316 8974
rect 5460 8945 5488 9862
rect 5264 8910 5316 8916
rect 5446 8936 5502 8945
rect 5276 8537 5304 8910
rect 5446 8871 5502 8880
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5262 8528 5318 8537
rect 5368 8498 5396 8774
rect 5262 8463 5318 8472
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 8090 5304 8230
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5276 6390 5304 7482
rect 5172 6384 5224 6390
rect 5078 6352 5134 6361
rect 5172 6326 5224 6332
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5078 6287 5134 6296
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 4146 5028 6190
rect 5092 5370 5120 6287
rect 5170 5944 5226 5953
rect 5170 5879 5226 5888
rect 5184 5710 5212 5879
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5368 5370 5396 8298
rect 5460 8090 5488 8871
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5644 6866 5672 12543
rect 5736 12238 5764 13942
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10062 5764 10406
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5736 8362 5764 8910
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5448 6656 5500 6662
rect 5736 6644 5764 7414
rect 5448 6598 5500 6604
rect 5552 6616 5764 6644
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4282 5396 4490
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4908 2774 4936 2994
rect 4816 2746 4936 2774
rect 4620 1828 4672 1834
rect 4620 1770 4672 1776
rect 4816 800 4844 2746
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 800 5212 2382
rect 5276 1630 5304 4014
rect 5460 2666 5488 6598
rect 5368 2638 5488 2666
rect 5368 1766 5396 2638
rect 5446 2544 5502 2553
rect 5446 2479 5448 2488
rect 5500 2479 5502 2488
rect 5448 2450 5500 2456
rect 5356 1760 5408 1766
rect 5356 1702 5408 1708
rect 5264 1624 5316 1630
rect 5264 1566 5316 1572
rect 5552 800 5580 6616
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 5409 5764 5646
rect 5722 5400 5778 5409
rect 5722 5335 5778 5344
rect 5630 4856 5686 4865
rect 5630 4791 5686 4800
rect 5644 4298 5672 4791
rect 5828 4706 5856 17070
rect 5920 16590 5948 17138
rect 6012 16726 6040 17274
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6012 15026 6040 15846
rect 6000 15020 6052 15026
rect 6104 15008 6132 17575
rect 6196 16266 6224 19207
rect 6288 17338 6316 22170
rect 7208 22114 7236 22578
rect 7104 22094 7156 22098
rect 7208 22094 7328 22114
rect 7104 22092 7328 22094
rect 7156 22086 7328 22092
rect 7156 22066 7236 22086
rect 7104 22034 7156 22040
rect 6550 21992 6606 22001
rect 6550 21927 6606 21936
rect 6736 21956 6788 21962
rect 6564 17796 6592 21927
rect 6736 21898 6788 21904
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 18698 6684 20742
rect 6748 20602 6776 21898
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6734 20496 6790 20505
rect 6840 20466 6868 21286
rect 7300 20466 7328 22086
rect 7484 21554 7512 24006
rect 7656 23792 7708 23798
rect 7656 23734 7708 23740
rect 7668 23186 7696 23734
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7668 22094 7696 22510
rect 7576 22066 7696 22094
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 6734 20431 6790 20440
rect 6828 20460 6880 20466
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6564 17768 6684 17796
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6472 16697 6500 17682
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6458 16688 6514 16697
rect 6458 16623 6514 16632
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6196 16238 6316 16266
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6196 15706 6224 16050
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6104 14980 6224 15008
rect 6000 14962 6052 14968
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6012 14074 6040 14486
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5920 11694 5948 13330
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12238 6040 12582
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5908 11688 5960 11694
rect 6000 11688 6052 11694
rect 5908 11630 5960 11636
rect 5998 11656 6000 11665
rect 6052 11656 6054 11665
rect 5998 11591 6054 11600
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 10266 5948 10610
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6012 10266 6040 10542
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5920 10062 5948 10202
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5906 8664 5962 8673
rect 5906 8599 5962 8608
rect 5920 8566 5948 8599
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7410 6040 8230
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5906 7304 5962 7313
rect 5906 7239 5962 7248
rect 5920 6798 5948 7239
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5736 4678 5856 4706
rect 5736 4434 5764 4678
rect 5736 4406 5856 4434
rect 5644 4270 5764 4298
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 4344 196 4396 202
rect 4344 138 4396 144
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5644 762 5672 4082
rect 5736 3670 5764 4270
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2514 5764 3130
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5828 2446 5856 4406
rect 5920 4146 5948 6734
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5906 4040 5962 4049
rect 5906 3975 5962 3984
rect 5920 3942 5948 3975
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 6012 3670 6040 7142
rect 6104 5234 6132 14826
rect 6196 12617 6224 14980
rect 6288 14906 6316 16238
rect 6380 16046 6408 16526
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6564 15008 6592 17546
rect 6656 16250 6684 17768
rect 6748 17082 6776 20431
rect 6828 20402 6880 20408
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19854 6960 20198
rect 7300 19854 7328 20402
rect 7378 20224 7434 20233
rect 7378 20159 7434 20168
rect 6920 19848 6972 19854
rect 7288 19848 7340 19854
rect 6972 19808 7144 19836
rect 6920 19790 6972 19796
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6840 17270 6868 17478
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6748 17054 6868 17082
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6748 16658 6776 16934
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6656 15570 6684 15982
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6840 15008 6868 17054
rect 6932 16522 6960 17478
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6932 15026 6960 15846
rect 7116 15450 7144 19808
rect 7288 19790 7340 19796
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 15586 7236 19654
rect 7300 19378 7328 19790
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7300 18834 7328 19314
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7300 18290 7328 18770
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7300 16046 7328 18226
rect 7392 16946 7420 20159
rect 7484 17678 7512 20742
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7392 16918 7512 16946
rect 7378 16824 7434 16833
rect 7378 16759 7434 16768
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7208 15570 7328 15586
rect 7208 15564 7340 15570
rect 7208 15558 7288 15564
rect 7288 15506 7340 15512
rect 7012 15428 7064 15434
rect 7116 15422 7236 15450
rect 7012 15370 7064 15376
rect 6472 14980 6592 15008
rect 6656 14980 6868 15008
rect 6920 15020 6972 15026
rect 6288 14878 6408 14906
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6288 14521 6316 14758
rect 6274 14512 6330 14521
rect 6274 14447 6330 14456
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6288 13530 6316 13874
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6380 12730 6408 14878
rect 6288 12702 6408 12730
rect 6182 12608 6238 12617
rect 6182 12543 6238 12552
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6196 10674 6224 10950
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4282 6132 5034
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6090 4040 6146 4049
rect 6090 3975 6146 3984
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5920 2446 5948 3334
rect 6104 3058 6132 3975
rect 6196 3074 6224 9590
rect 6288 6730 6316 12702
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 9110 6408 12582
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6380 5658 6408 8502
rect 6472 7041 6500 14980
rect 6550 14920 6606 14929
rect 6550 14855 6552 14864
rect 6604 14855 6606 14864
rect 6552 14826 6604 14832
rect 6550 14648 6606 14657
rect 6550 14583 6606 14592
rect 6564 14278 6592 14583
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 14074 6592 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6656 12730 6684 14980
rect 6920 14962 6972 14968
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13326 6776 14214
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6840 12782 6868 14826
rect 7024 14618 7052 15370
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 14498 7144 15302
rect 7208 15065 7236 15422
rect 7194 15056 7250 15065
rect 7194 14991 7250 15000
rect 7392 14550 7420 16759
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7024 14470 7144 14498
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 6932 13841 6960 14418
rect 6918 13832 6974 13841
rect 6918 13767 6974 13776
rect 6564 12702 6684 12730
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6564 12646 6592 12702
rect 6552 12640 6604 12646
rect 6644 12640 6696 12646
rect 6552 12582 6604 12588
rect 6642 12608 6644 12617
rect 6696 12608 6698 12617
rect 6642 12543 6698 12552
rect 6656 11830 6684 12543
rect 6840 11830 6868 12718
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11529 6960 11562
rect 6918 11520 6974 11529
rect 6918 11455 6974 11464
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 6564 6934 6592 11290
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10169 6684 11086
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6748 10656 6776 10746
rect 6920 10668 6972 10674
rect 6748 10628 6920 10656
rect 6920 10610 6972 10616
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6642 10160 6698 10169
rect 6642 10095 6698 10104
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6656 8566 6684 9114
rect 6748 8906 6776 10474
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6826 8936 6882 8945
rect 6736 8900 6788 8906
rect 6826 8871 6882 8880
rect 6736 8842 6788 8848
rect 6840 8634 6868 8871
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 7449 6868 7482
rect 6826 7440 6882 7449
rect 6826 7375 6882 7384
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 7041 6684 7142
rect 6642 7032 6698 7041
rect 6642 6967 6698 6976
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6288 5630 6408 5658
rect 6288 3194 6316 5630
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6092 3052 6144 3058
rect 6196 3046 6316 3074
rect 6092 2994 6144 3000
rect 6184 2984 6236 2990
rect 6182 2952 6184 2961
rect 6236 2952 6238 2961
rect 6182 2887 6238 2896
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 5828 870 5948 898
rect 5828 762 5856 870
rect 5920 800 5948 870
rect 5644 734 5856 762
rect 5906 0 5962 800
rect 6196 134 6224 2887
rect 6288 800 6316 3046
rect 6380 2417 6408 5510
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6366 2408 6422 2417
rect 6366 2343 6422 2352
rect 6472 1222 6500 3878
rect 6564 2938 6592 6734
rect 6656 4486 6684 6967
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6748 6118 6776 6190
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6642 3632 6698 3641
rect 6642 3567 6698 3576
rect 6656 3194 6684 3567
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6748 3074 6776 6054
rect 6840 5914 6868 6054
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6840 3194 6868 3470
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6748 3046 6868 3074
rect 6932 3058 6960 10406
rect 7024 10305 7052 14470
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7116 12442 7144 14282
rect 7392 13138 7420 14282
rect 7484 13258 7512 16918
rect 7576 15201 7604 22066
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7562 15192 7618 15201
rect 7562 15127 7618 15136
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7576 14618 7604 14758
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7668 14346 7696 20878
rect 7760 20058 7788 32846
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8864 28762 8892 38898
rect 9048 32570 9076 45358
rect 9128 35692 9180 35698
rect 9128 35634 9180 35640
rect 9036 32564 9088 32570
rect 9036 32506 9088 32512
rect 8852 28756 8904 28762
rect 8852 28698 8904 28704
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 8680 28082 8708 28494
rect 8668 28076 8720 28082
rect 8588 28036 8668 28064
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 7840 23180 7892 23186
rect 8404 23168 8432 23462
rect 8496 23322 8524 26318
rect 8588 24818 8616 28036
rect 8668 28018 8720 28024
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8956 26586 8984 27950
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8944 25696 8996 25702
rect 8944 25638 8996 25644
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 8956 25498 8984 25638
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8942 24712 8998 24721
rect 8942 24647 8998 24656
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8404 23140 8524 23168
rect 7840 23122 7892 23128
rect 7852 22642 7880 23122
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 8496 22506 8524 23140
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7852 20942 7880 22374
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8220 21876 8248 21966
rect 8220 21848 8340 21876
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8312 21672 8340 21848
rect 8220 21644 8340 21672
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 8220 20856 8248 21644
rect 8220 20828 8340 20856
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8116 20528 8168 20534
rect 8114 20496 8116 20505
rect 8168 20496 8170 20505
rect 8114 20431 8170 20440
rect 7748 20052 7800 20058
rect 7932 20052 7984 20058
rect 7748 19994 7800 20000
rect 7852 20012 7932 20040
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7760 17746 7788 19858
rect 7852 19446 7880 20012
rect 7932 19994 7984 20000
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 19446 8340 20828
rect 8390 20360 8446 20369
rect 8390 20295 8446 20304
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 7932 19304 7984 19310
rect 7852 19264 7932 19292
rect 7852 17882 7880 19264
rect 8312 19258 8340 19382
rect 7932 19246 7984 19252
rect 8128 19230 8340 19258
rect 8128 18834 8156 19230
rect 8208 19168 8260 19174
rect 8404 19122 8432 20295
rect 8496 19922 8524 22442
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8680 21622 8708 21830
rect 8864 21690 8892 22510
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8668 21616 8720 21622
rect 8668 21558 8720 21564
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8588 19514 8616 20198
rect 8666 20088 8722 20097
rect 8956 20040 8984 24647
rect 9048 20244 9076 25638
rect 9140 23866 9168 35634
rect 9324 33114 9352 45902
rect 9496 45554 9548 45558
rect 9600 45554 9628 47126
rect 9772 47048 9824 47054
rect 9772 46990 9824 46996
rect 9784 46170 9812 46990
rect 9772 46164 9824 46170
rect 9772 46106 9824 46112
rect 10152 46034 10180 48486
rect 10508 47456 10560 47462
rect 10508 47398 10560 47404
rect 10324 47252 10376 47258
rect 10324 47194 10376 47200
rect 10140 46028 10192 46034
rect 10140 45970 10192 45976
rect 9496 45552 9628 45554
rect 9548 45526 9628 45552
rect 9496 45494 9548 45500
rect 10152 45082 10180 45970
rect 10140 45076 10192 45082
rect 10140 45018 10192 45024
rect 10232 44396 10284 44402
rect 10232 44338 10284 44344
rect 10244 43994 10272 44338
rect 10232 43988 10284 43994
rect 10232 43930 10284 43936
rect 10336 43790 10364 47194
rect 10520 44878 10548 47398
rect 10796 46034 10824 51954
rect 10784 46028 10836 46034
rect 10784 45970 10836 45976
rect 10796 45626 10824 45970
rect 10784 45620 10836 45626
rect 10784 45562 10836 45568
rect 10980 45422 11008 56222
rect 12070 56200 12126 57000
rect 13450 56200 13506 57000
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 16316 56222 16528 56250
rect 11060 54120 11112 54126
rect 11060 54062 11112 54068
rect 11072 50726 11100 54062
rect 11060 50720 11112 50726
rect 11060 50662 11112 50668
rect 11072 48822 11100 50662
rect 11428 48884 11480 48890
rect 11428 48826 11480 48832
rect 11060 48816 11112 48822
rect 11060 48758 11112 48764
rect 11072 47258 11100 48758
rect 11440 48142 11468 48826
rect 11428 48136 11480 48142
rect 11428 48078 11480 48084
rect 11428 48000 11480 48006
rect 11428 47942 11480 47948
rect 11060 47252 11112 47258
rect 11060 47194 11112 47200
rect 11072 47054 11100 47194
rect 11060 47048 11112 47054
rect 11060 46990 11112 46996
rect 11072 45554 11100 46990
rect 11440 46646 11468 47942
rect 11428 46640 11480 46646
rect 11428 46582 11480 46588
rect 12084 46034 12112 56200
rect 13464 54194 13492 56200
rect 14844 54194 14872 56200
rect 16224 56114 16252 56200
rect 16316 56114 16344 56222
rect 16224 56086 16344 56114
rect 16500 54210 16528 56222
rect 17590 56200 17646 57000
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 21730 56200 21786 57000
rect 22848 56222 23060 56250
rect 16500 54194 16620 54210
rect 17604 54194 17632 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18984 54330 19012 56200
rect 18972 54324 19024 54330
rect 18972 54266 19024 54272
rect 13452 54188 13504 54194
rect 13452 54130 13504 54136
rect 14832 54188 14884 54194
rect 16500 54188 16632 54194
rect 16500 54182 16580 54188
rect 14832 54130 14884 54136
rect 16580 54130 16632 54136
rect 17592 54188 17644 54194
rect 17592 54130 17644 54136
rect 18984 54126 19012 54266
rect 18972 54120 19024 54126
rect 18972 54062 19024 54068
rect 16764 54052 16816 54058
rect 16764 53994 16816 54000
rect 13544 53984 13596 53990
rect 13544 53926 13596 53932
rect 14924 53984 14976 53990
rect 14924 53926 14976 53932
rect 15660 53984 15712 53990
rect 15660 53926 15712 53932
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12164 47048 12216 47054
rect 12164 46990 12216 46996
rect 12072 46028 12124 46034
rect 12072 45970 12124 45976
rect 12176 45626 12204 46990
rect 13556 46510 13584 53926
rect 14464 48000 14516 48006
rect 14464 47942 14516 47948
rect 14476 46986 14504 47942
rect 14648 47456 14700 47462
rect 14648 47398 14700 47404
rect 14280 46980 14332 46986
rect 14280 46922 14332 46928
rect 14464 46980 14516 46986
rect 14464 46922 14516 46928
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 14292 46034 14320 46922
rect 14660 46646 14688 47398
rect 14936 47122 14964 53926
rect 14924 47116 14976 47122
rect 14924 47058 14976 47064
rect 14648 46640 14700 46646
rect 14648 46582 14700 46588
rect 15672 46510 15700 53926
rect 16212 53100 16264 53106
rect 16212 53042 16264 53048
rect 15660 46504 15712 46510
rect 15660 46446 15712 46452
rect 14280 46028 14332 46034
rect 14280 45970 14332 45976
rect 12164 45620 12216 45626
rect 12164 45562 12216 45568
rect 11072 45526 11192 45554
rect 11164 45490 11192 45526
rect 11152 45484 11204 45490
rect 11152 45426 11204 45432
rect 10968 45416 11020 45422
rect 10968 45358 11020 45364
rect 11796 45280 11848 45286
rect 11796 45222 11848 45228
rect 11520 44940 11572 44946
rect 11520 44882 11572 44888
rect 10508 44872 10560 44878
rect 10508 44814 10560 44820
rect 10876 44872 10928 44878
rect 10876 44814 10928 44820
rect 10520 44198 10548 44814
rect 10888 44538 10916 44814
rect 10876 44532 10928 44538
rect 10876 44474 10928 44480
rect 11532 44334 11560 44882
rect 11520 44328 11572 44334
rect 11520 44270 11572 44276
rect 10508 44192 10560 44198
rect 10508 44134 10560 44140
rect 9956 43784 10008 43790
rect 9956 43726 10008 43732
rect 10324 43784 10376 43790
rect 10324 43726 10376 43732
rect 9968 42566 9996 43726
rect 11532 42770 11560 44270
rect 11520 42764 11572 42770
rect 11520 42706 11572 42712
rect 11532 42566 11560 42706
rect 9956 42560 10008 42566
rect 9956 42502 10008 42508
rect 11520 42560 11572 42566
rect 11520 42502 11572 42508
rect 11244 39432 11296 39438
rect 11244 39374 11296 39380
rect 11256 38010 11284 39374
rect 11244 38004 11296 38010
rect 11244 37946 11296 37952
rect 11152 37868 11204 37874
rect 11152 37810 11204 37816
rect 11164 35630 11192 37810
rect 11532 35894 11560 42502
rect 11808 37874 11836 45222
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 14372 44260 14424 44266
rect 14372 44202 14424 44208
rect 11980 44192 12032 44198
rect 11980 44134 12032 44140
rect 11992 43722 12020 44134
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 11980 43716 12032 43722
rect 11980 43658 12032 43664
rect 11888 42900 11940 42906
rect 11888 42842 11940 42848
rect 11900 39642 11928 42842
rect 11992 42770 12020 43658
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 11980 42764 12032 42770
rect 11980 42706 12032 42712
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 14384 41414 14412 44202
rect 15936 42764 15988 42770
rect 15936 42706 15988 42712
rect 14108 41386 14412 41414
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 11888 39636 11940 39642
rect 11888 39578 11940 39584
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 11796 37868 11848 37874
rect 11796 37810 11848 37816
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 11532 35866 11652 35894
rect 11532 35834 11560 35866
rect 11520 35828 11572 35834
rect 11520 35770 11572 35776
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 11152 35624 11204 35630
rect 11152 35566 11204 35572
rect 9692 34202 9720 35566
rect 11624 35494 11652 35866
rect 11704 35760 11756 35766
rect 11704 35702 11756 35708
rect 11612 35488 11664 35494
rect 11612 35430 11664 35436
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 11624 34066 11652 35430
rect 11612 34060 11664 34066
rect 11612 34002 11664 34008
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9220 32428 9272 32434
rect 9220 32370 9272 32376
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 9140 22137 9168 22646
rect 9126 22128 9182 22137
rect 9126 22063 9182 22072
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9140 20398 9168 20810
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9048 20216 9168 20244
rect 8666 20023 8722 20032
rect 8680 19825 8708 20023
rect 8772 20012 8984 20040
rect 8666 19816 8722 19825
rect 8666 19751 8722 19760
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8260 19116 8432 19122
rect 8208 19110 8432 19116
rect 8220 19094 8432 19110
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8404 18358 8432 18770
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 16794 7788 17682
rect 8496 17610 8524 19450
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8588 18766 8616 19178
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8588 18358 8616 18702
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 16998 8340 17070
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7930 16552 7986 16561
rect 7930 16487 7986 16496
rect 7944 16454 7972 16487
rect 7932 16448 7984 16454
rect 8220 16436 8248 16934
rect 8300 16720 8352 16726
rect 8298 16688 8300 16697
rect 8352 16688 8354 16697
rect 8298 16623 8354 16632
rect 8588 16522 8616 18294
rect 8576 16516 8628 16522
rect 8576 16458 8628 16464
rect 8484 16448 8536 16454
rect 8220 16408 8340 16436
rect 7932 16390 7984 16396
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7760 16114 7788 16186
rect 8312 16182 8340 16408
rect 8482 16416 8484 16425
rect 8536 16416 8538 16425
rect 8482 16351 8538 16360
rect 8588 16266 8616 16458
rect 8496 16238 8616 16266
rect 8496 16182 8524 16238
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7852 15026 7880 15914
rect 7944 15473 7972 15914
rect 8128 15473 8156 16118
rect 8220 15966 8432 15994
rect 7930 15464 7986 15473
rect 7930 15399 7986 15408
rect 8114 15464 8170 15473
rect 8114 15399 8170 15408
rect 8220 15348 8248 15966
rect 8404 15910 8432 15966
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8390 15600 8446 15609
rect 8390 15535 8446 15544
rect 8220 15320 8340 15348
rect 8404 15337 8432 15535
rect 8588 15502 8616 16238
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7930 15056 7986 15065
rect 7840 15020 7892 15026
rect 7930 14991 7986 15000
rect 7840 14962 7892 14968
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7760 14278 7788 14826
rect 7944 14328 7972 14991
rect 7852 14300 7972 14328
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 14006 7788 14214
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7852 13954 7880 14300
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7852 13926 8156 13954
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7748 13524 7800 13530
rect 7932 13524 7984 13530
rect 7800 13484 7932 13512
rect 7748 13466 7800 13472
rect 7932 13466 7984 13472
rect 8036 13326 8064 13738
rect 8128 13326 8156 13926
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7748 13184 7800 13190
rect 7392 13110 7696 13138
rect 7932 13184 7984 13190
rect 7800 13144 7932 13172
rect 7748 13126 7800 13132
rect 7932 13126 7984 13132
rect 7668 12782 7696 13110
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7576 12481 7604 12718
rect 7760 12646 7788 12922
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7562 12472 7618 12481
rect 7104 12436 7156 12442
rect 7562 12407 7618 12416
rect 7104 12378 7156 12384
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7010 10296 7066 10305
rect 7010 10231 7066 10240
rect 7116 10180 7144 11494
rect 7668 11354 7696 11630
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7470 11248 7526 11257
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7380 11212 7432 11218
rect 7470 11183 7526 11192
rect 7380 11154 7432 11160
rect 7300 10742 7328 11154
rect 7288 10736 7340 10742
rect 7286 10704 7288 10713
rect 7340 10704 7342 10713
rect 7286 10639 7342 10648
rect 7024 10152 7144 10180
rect 7024 7970 7052 10152
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 8090 7144 9930
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9058 7236 9862
rect 7300 9654 7328 9998
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7392 9602 7420 11154
rect 7484 10742 7512 11183
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7760 10470 7788 12310
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 12102 8064 12174
rect 8220 12170 8248 12650
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8128 11694 8156 11766
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8312 11506 8340 15320
rect 8390 15328 8446 15337
rect 8390 15263 8446 15272
rect 8496 15178 8524 15370
rect 8404 15150 8524 15178
rect 8404 15094 8432 15150
rect 8588 15094 8616 15438
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8404 13870 8432 15030
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8220 11478 8340 11506
rect 8220 11218 8248 11478
rect 8298 11384 8354 11393
rect 8404 11354 8432 13670
rect 8588 12850 8616 13670
rect 8680 12986 8708 18702
rect 8772 15706 8800 20012
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 16454 8892 19654
rect 8956 17338 8984 19722
rect 9048 19553 9076 19858
rect 9034 19544 9090 19553
rect 9034 19479 9090 19488
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8772 15502 8800 15642
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8956 15314 8984 17138
rect 9048 16289 9076 18566
rect 9140 17746 9168 20216
rect 9232 19786 9260 32370
rect 9784 32026 9812 33934
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 10508 31884 10560 31890
rect 10508 31826 10560 31832
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 9692 30326 9720 31758
rect 10324 31204 10376 31210
rect 10324 31146 10376 31152
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9680 30320 9732 30326
rect 9680 30262 9732 30268
rect 9784 29238 9812 31078
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10152 29481 10180 30670
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10138 29472 10194 29481
rect 10138 29407 10194 29416
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9416 28558 9444 29038
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9312 27328 9364 27334
rect 9310 27296 9312 27305
rect 9364 27296 9366 27305
rect 9310 27231 9366 27240
rect 9324 26994 9352 27231
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9416 26586 9444 26930
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9324 19242 9352 19654
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18057 9260 18566
rect 9416 18442 9444 23122
rect 9508 19514 9536 26250
rect 9692 25974 9720 26726
rect 9968 26234 9996 28358
rect 9968 26206 10088 26234
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9680 25220 9732 25226
rect 9680 25162 9732 25168
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9600 24206 9628 24890
rect 9692 24596 9720 25162
rect 9864 24608 9916 24614
rect 9692 24568 9864 24596
rect 9864 24550 9916 24556
rect 10060 24410 10088 26206
rect 10152 25498 10180 29407
rect 10244 28626 10272 30194
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 10244 28218 10272 28562
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10336 27674 10364 31146
rect 10520 30258 10548 31826
rect 11152 31816 11204 31822
rect 11152 31758 11204 31764
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 11072 29714 11100 30534
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10692 28688 10744 28694
rect 10692 28630 10744 28636
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10232 27056 10284 27062
rect 10232 26998 10284 27004
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 9680 23656 9732 23662
rect 9600 23616 9680 23644
rect 9600 22030 9628 23616
rect 9680 23598 9732 23604
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9692 21690 9720 22986
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9600 18902 9628 20266
rect 9692 20058 9720 20946
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9324 18414 9444 18442
rect 9692 18426 9720 19994
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9680 18420 9732 18426
rect 9218 18048 9274 18057
rect 9218 17983 9274 17992
rect 9324 17882 9352 18414
rect 9680 18362 9732 18368
rect 9678 18320 9734 18329
rect 9678 18255 9734 18264
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9034 16280 9090 16289
rect 9034 16215 9090 16224
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8864 15286 8984 15314
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8772 13802 8800 14758
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8298 11319 8354 11328
rect 8392 11348 8444 11354
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10470 8064 10610
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7760 9674 7788 10134
rect 7944 10010 7972 10406
rect 7668 9654 7788 9674
rect 7656 9648 7788 9654
rect 7392 9574 7512 9602
rect 7708 9646 7788 9648
rect 7852 9982 7972 10010
rect 7656 9590 7708 9596
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7208 9030 7328 9058
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7208 8634 7236 8910
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7024 7942 7144 7970
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 7177 7052 7278
rect 7010 7168 7066 7177
rect 7010 7103 7066 7112
rect 7116 6905 7144 7942
rect 7300 7857 7328 9030
rect 7392 8362 7420 9386
rect 7484 8634 7512 9574
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7576 8566 7604 9454
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7668 8498 7696 9318
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7484 8090 7512 8434
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7286 7848 7342 7857
rect 7286 7783 7342 7792
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7102 6896 7158 6905
rect 7102 6831 7158 6840
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 4146 7052 6122
rect 7116 5234 7144 6598
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5914 7236 6258
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7288 5840 7340 5846
rect 7208 5788 7288 5794
rect 7208 5782 7340 5788
rect 7208 5766 7328 5782
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6564 2910 6684 2938
rect 6460 1216 6512 1222
rect 6460 1158 6512 1164
rect 6656 800 6684 2910
rect 6840 1465 6868 3046
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6826 1456 6882 1465
rect 6826 1391 6882 1400
rect 7024 800 7052 3674
rect 7116 3670 7144 4218
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7208 1970 7236 5766
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 7300 2378 7328 5607
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 3738 7420 5306
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7484 3505 7512 7346
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 5710 7604 7142
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7668 5896 7696 6326
rect 7760 6066 7788 8570
rect 7852 6372 7880 9982
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8312 9674 8340 11319
rect 8392 11290 8444 11296
rect 8496 11218 8524 12718
rect 8772 12714 8800 13194
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8758 12472 8814 12481
rect 8758 12407 8814 12416
rect 8772 12102 8800 12407
rect 8864 12238 8892 15286
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8956 14958 8984 15098
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8956 13326 8984 14418
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8588 11150 8616 12038
rect 8668 11688 8720 11694
rect 8772 11676 8800 12038
rect 8720 11648 8800 11676
rect 8668 11630 8720 11636
rect 8956 11626 8984 13126
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8404 10266 8432 11086
rect 8482 10704 8538 10713
rect 8482 10639 8538 10648
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8496 10130 8524 10639
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8220 9353 8248 9658
rect 8312 9646 8432 9674
rect 8206 9344 8262 9353
rect 8206 9279 8262 9288
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8312 8634 8340 8910
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8404 8430 8432 9646
rect 8482 9208 8538 9217
rect 8482 9143 8538 9152
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8496 8242 8524 9143
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8566 8616 8774
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8404 8214 8524 8242
rect 7930 8120 7986 8129
rect 7930 8055 7986 8064
rect 7944 8022 7972 8055
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7852 6344 7972 6372
rect 7760 6038 7880 6066
rect 7668 5868 7788 5896
rect 7654 5808 7710 5817
rect 7760 5778 7788 5868
rect 7654 5743 7656 5752
rect 7708 5743 7710 5752
rect 7748 5772 7800 5778
rect 7656 5714 7708 5720
rect 7748 5714 7800 5720
rect 7564 5704 7616 5710
rect 7852 5658 7880 6038
rect 7944 5681 7972 6344
rect 7564 5646 7616 5652
rect 7760 5630 7880 5658
rect 7930 5672 7986 5681
rect 7562 5536 7618 5545
rect 7562 5471 7618 5480
rect 7470 3496 7526 3505
rect 7470 3431 7526 3440
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 7392 800 7420 3062
rect 7484 882 7512 3334
rect 7576 2106 7604 5471
rect 7654 5400 7710 5409
rect 7654 5335 7656 5344
rect 7708 5335 7710 5344
rect 7656 5306 7708 5312
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7668 4826 7696 5199
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7668 4282 7696 4422
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7760 4026 7788 5630
rect 7930 5607 7986 5616
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 8312 4729 8340 7822
rect 8298 4720 8354 4729
rect 8404 4706 8432 8214
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 4826 8524 7686
rect 8574 7576 8630 7585
rect 8574 7511 8630 7520
rect 8588 7478 8616 7511
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8574 6896 8630 6905
rect 8574 6831 8630 6840
rect 8588 6633 8616 6831
rect 8574 6624 8630 6633
rect 8574 6559 8630 6568
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8404 4678 8524 4706
rect 8298 4655 8354 4664
rect 8496 4622 8524 4678
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8404 4321 8432 4558
rect 8482 4448 8538 4457
rect 8482 4383 8538 4392
rect 8390 4312 8446 4321
rect 8390 4247 8446 4256
rect 7668 3998 7788 4026
rect 7668 3369 7696 3998
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7654 3360 7710 3369
rect 7654 3295 7710 3304
rect 7654 3224 7710 3233
rect 7654 3159 7710 3168
rect 7668 3126 7696 3159
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7760 2394 7788 3878
rect 7930 3632 7986 3641
rect 7930 3567 7986 3576
rect 7944 3534 7972 3567
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8312 3058 8340 3334
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7668 2366 7788 2394
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7668 950 7696 2366
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7656 944 7708 950
rect 7656 886 7708 892
rect 7472 876 7524 882
rect 7472 818 7524 824
rect 7760 800 7788 2246
rect 7852 1018 7880 2926
rect 8300 2848 8352 2854
rect 8298 2816 8300 2825
rect 8352 2816 8354 2825
rect 8298 2751 8354 2760
rect 8496 2774 8524 4383
rect 8588 2990 8616 6054
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 7932 1352 7984 1358
rect 7930 1320 7932 1329
rect 7984 1320 7986 1329
rect 7930 1255 7986 1264
rect 7840 1012 7892 1018
rect 7840 954 7892 960
rect 8128 800 8156 2042
rect 8312 1086 8340 2751
rect 8496 2746 8616 2774
rect 8390 2680 8446 2689
rect 8390 2615 8446 2624
rect 8404 2145 8432 2615
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8390 2136 8446 2145
rect 8390 2071 8446 2080
rect 8300 1080 8352 1086
rect 8300 1022 8352 1028
rect 8496 800 8524 2450
rect 8588 1170 8616 2746
rect 8680 1290 8708 10202
rect 8772 9518 8800 11494
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8864 10810 8892 11018
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8772 8430 8800 9454
rect 8956 9178 8984 11018
rect 9048 10146 9076 15642
rect 9140 13870 9168 17206
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9232 13530 9260 16594
rect 9416 15638 9444 17070
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 15706 9536 16526
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9404 15632 9456 15638
rect 9404 15574 9456 15580
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9324 14482 9352 15098
rect 9508 14482 9536 15370
rect 9600 15162 9628 17546
rect 9692 17542 9720 18255
rect 9784 17785 9812 19382
rect 9968 18465 9996 21966
rect 9954 18456 10010 18465
rect 9954 18391 10010 18400
rect 9968 18358 9996 18391
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9770 17776 9826 17785
rect 9770 17711 9826 17720
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9954 17504 10010 17513
rect 9954 17439 10010 17448
rect 9968 17338 9996 17439
rect 10060 17338 10088 23802
rect 10152 23662 10180 25094
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 10152 20534 10180 22646
rect 10244 21894 10272 26998
rect 10324 26512 10376 26518
rect 10322 26480 10324 26489
rect 10376 26480 10378 26489
rect 10322 26415 10378 26424
rect 10324 25832 10376 25838
rect 10324 25774 10376 25780
rect 10336 23866 10364 25774
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10336 21146 10364 23666
rect 10428 21690 10456 28358
rect 10520 26994 10548 28426
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10704 26874 10732 28630
rect 10888 27538 10916 29582
rect 11164 29034 11192 31758
rect 11244 31340 11296 31346
rect 11244 31282 11296 31288
rect 11256 30938 11284 31282
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 11716 30394 11744 35702
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13912 32020 13964 32026
rect 13912 31962 13964 31968
rect 12072 31952 12124 31958
rect 12072 31894 12124 31900
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 11520 29572 11572 29578
rect 11520 29514 11572 29520
rect 11716 29560 11744 30330
rect 11808 30326 11836 30670
rect 11796 30320 11848 30326
rect 11796 30262 11848 30268
rect 11796 29572 11848 29578
rect 11716 29532 11796 29560
rect 11532 29306 11560 29514
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11716 29238 11744 29532
rect 11796 29514 11848 29520
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11152 29028 11204 29034
rect 11152 28970 11204 28976
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 11072 28082 11100 28494
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 10966 27976 11022 27985
rect 10966 27911 11022 27920
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 10980 26926 11008 27911
rect 11164 26926 11192 28970
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11336 28484 11388 28490
rect 11336 28426 11388 28432
rect 11348 27130 11376 28426
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 10520 26846 10732 26874
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 10520 25922 10548 26846
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10612 26081 10640 26386
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10598 26072 10654 26081
rect 10598 26007 10654 26016
rect 10520 25894 10732 25922
rect 10704 25838 10732 25894
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10508 25424 10560 25430
rect 10508 25366 10560 25372
rect 10520 24954 10548 25366
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10508 24064 10560 24070
rect 10508 24006 10560 24012
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10140 20528 10192 20534
rect 10140 20470 10192 20476
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10138 17776 10194 17785
rect 10138 17711 10194 17720
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9692 16522 9720 16934
rect 9784 16697 9812 16934
rect 9770 16688 9826 16697
rect 9770 16623 9826 16632
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14550 9628 14962
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9784 14414 9812 15982
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 14278 9812 14350
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9140 10266 9168 13262
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9232 11626 9260 11834
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9324 10742 9352 13330
rect 9416 12986 9444 14010
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9416 12850 9444 12922
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9416 11694 9444 12786
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9508 11354 9536 14010
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 11898 9628 13738
rect 9784 13394 9812 13806
rect 9876 13530 9904 17206
rect 10152 16969 10180 17711
rect 10336 17134 10364 18362
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10138 16960 10194 16969
rect 10138 16895 10194 16904
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 9954 16280 10010 16289
rect 9954 16215 9956 16224
rect 10008 16215 10010 16224
rect 9956 16186 10008 16192
rect 9968 15094 9996 16186
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 10060 14074 10088 16390
rect 10152 16182 10180 16390
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10152 15910 10180 16118
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10152 15366 10180 15574
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10244 13802 10272 13942
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13569 9996 13670
rect 9954 13560 10010 13569
rect 9864 13524 9916 13530
rect 9954 13495 10010 13504
rect 9864 13466 9916 13472
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9692 12434 9720 13330
rect 9784 13190 9812 13330
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9770 13016 9826 13025
rect 9770 12951 9826 12960
rect 9784 12918 9812 12951
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10152 12481 10180 12854
rect 10138 12472 10194 12481
rect 9864 12436 9916 12442
rect 9692 12406 9812 12434
rect 9784 12238 9812 12406
rect 10138 12407 10194 12416
rect 9864 12378 9916 12384
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 12073 9720 12106
rect 9678 12064 9734 12073
rect 9678 11999 9734 12008
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9876 11150 9904 12378
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 10060 11898 10088 12310
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10152 10742 10180 12407
rect 10336 11529 10364 15030
rect 10428 11744 10456 19450
rect 10520 18426 10548 24006
rect 10612 22166 10640 25434
rect 10796 25226 10824 25842
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 10796 24886 10824 25162
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10704 23186 10732 24550
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10796 23050 10824 24822
rect 10888 24614 10916 26318
rect 11336 26036 11388 26042
rect 11336 25978 11388 25984
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10980 25362 11008 25910
rect 11348 25906 11376 25978
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10796 22710 10824 22986
rect 10888 22982 10916 24210
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10704 22030 10732 22374
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10888 21842 10916 22918
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 21978 11008 22510
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22094 11100 22374
rect 11072 22066 11192 22094
rect 10980 21950 11100 21978
rect 10612 20602 10640 21830
rect 10796 21434 10824 21830
rect 10888 21814 11008 21842
rect 10980 21486 11008 21814
rect 11072 21554 11100 21950
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10968 21480 11020 21486
rect 10796 21418 10916 21434
rect 10968 21422 11020 21428
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10796 21412 10928 21418
rect 10796 21406 10876 21412
rect 10704 21146 10732 21354
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10612 18834 10640 19110
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 13530 10548 14214
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10520 11937 10548 12922
rect 10612 12442 10640 18770
rect 10704 16250 10732 20742
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10796 16182 10824 21406
rect 10876 21354 10928 21360
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20466 11100 20878
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11164 20040 11192 22066
rect 11256 21418 11284 24142
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11256 21010 11284 21354
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11072 20012 11192 20040
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10888 15201 10916 19110
rect 11072 18766 11100 20012
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10968 17876 11020 17882
rect 11072 17864 11100 18566
rect 11020 17836 11100 17864
rect 10968 17818 11020 17824
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16182 11100 16662
rect 11164 16658 11192 19858
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11348 18986 11376 19654
rect 11440 19378 11468 28562
rect 11716 28506 11744 29174
rect 11900 29170 11928 29446
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11716 28490 11836 28506
rect 11716 28484 11848 28490
rect 11716 28478 11796 28484
rect 11716 28218 11744 28478
rect 11796 28426 11848 28432
rect 11704 28212 11756 28218
rect 11704 28154 11756 28160
rect 11716 27674 11744 28154
rect 11704 27668 11756 27674
rect 11704 27610 11756 27616
rect 11716 27402 11744 27610
rect 11704 27396 11756 27402
rect 11704 27338 11756 27344
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11624 26450 11652 27270
rect 12084 26994 12112 31894
rect 12624 31884 12676 31890
rect 12624 31826 12676 31832
rect 12636 30190 12664 31826
rect 13544 31748 13596 31754
rect 13544 31690 13596 31696
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12716 30660 12768 30666
rect 12716 30602 12768 30608
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12452 27130 12480 27950
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 11612 26444 11664 26450
rect 11612 26386 11664 26392
rect 11520 26308 11572 26314
rect 11520 26250 11572 26256
rect 11532 24274 11560 26250
rect 11624 25906 11652 26386
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11716 24818 11744 25638
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11348 18958 11468 18986
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11348 18630 11376 18838
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11440 18442 11468 18958
rect 11348 18414 11468 18442
rect 11532 18426 11560 21014
rect 11520 18420 11572 18426
rect 11348 17882 11376 18414
rect 11520 18362 11572 18368
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11336 17876 11388 17882
rect 11256 17836 11336 17864
rect 11256 17610 11284 17836
rect 11336 17818 11388 17824
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11348 17270 11376 17682
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11242 15872 11298 15881
rect 11242 15807 11298 15816
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10874 15192 10930 15201
rect 10874 15127 10930 15136
rect 10874 14104 10930 14113
rect 10874 14039 10876 14048
rect 10928 14039 10930 14048
rect 10876 14010 10928 14016
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10704 13802 10732 13874
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10600 12436 10652 12442
rect 10796 12434 10824 13738
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10600 12378 10652 12384
rect 10704 12406 10824 12434
rect 10704 12170 10732 12406
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10506 11928 10562 11937
rect 10506 11863 10562 11872
rect 10508 11756 10560 11762
rect 10428 11716 10508 11744
rect 10428 11558 10456 11716
rect 10508 11698 10560 11704
rect 10416 11552 10468 11558
rect 10322 11520 10378 11529
rect 10416 11494 10468 11500
rect 10322 11455 10378 11464
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9312 10600 9364 10606
rect 9364 10560 9444 10588
rect 9312 10542 9364 10548
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9048 10118 9352 10146
rect 9416 10130 9444 10560
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9324 10010 9352 10118
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9048 9722 9076 9998
rect 9324 9994 9536 10010
rect 9324 9988 9548 9994
rect 9324 9982 9496 9988
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 9178 9168 9454
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8850 9072 8906 9081
rect 8850 9007 8852 9016
rect 8904 9007 8906 9016
rect 8852 8978 8904 8984
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8772 7342 8800 8366
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8942 8120 8998 8129
rect 8942 8055 8998 8064
rect 9036 8084 9088 8090
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8864 6798 8892 7686
rect 8956 7002 8984 8055
rect 9036 8026 9088 8032
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8772 6458 8800 6734
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5710 8984 6054
rect 8944 5704 8996 5710
rect 8758 5672 8814 5681
rect 8944 5646 8996 5652
rect 8758 5607 8814 5616
rect 8772 4214 8800 5607
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8864 4321 8892 4966
rect 8850 4312 8906 4321
rect 8850 4247 8906 4256
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8956 4146 8984 4966
rect 9048 4826 9076 8026
rect 9140 7886 9168 8026
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9232 6866 9260 8230
rect 9324 7886 9352 9982
rect 9496 9930 9548 9936
rect 9588 9920 9640 9926
rect 9586 9888 9588 9897
rect 9640 9888 9642 9897
rect 9586 9823 9642 9832
rect 9404 9648 9456 9654
rect 9456 9608 9536 9636
rect 9404 9590 9456 9596
rect 9508 8974 9536 9608
rect 9784 9518 9812 10066
rect 10152 9994 10180 10678
rect 10336 10470 10364 11154
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 10152 9450 10180 9930
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 7954 9720 8774
rect 10152 8498 10180 9386
rect 10244 9110 10272 10406
rect 10428 9761 10456 10950
rect 10414 9752 10470 9761
rect 10414 9687 10470 9696
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10428 9450 10456 9522
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10520 8974 10548 11018
rect 10612 10849 10640 12106
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10704 11014 10732 11834
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10598 10840 10654 10849
rect 10598 10775 10654 10784
rect 10612 10282 10640 10775
rect 10612 10266 10732 10282
rect 10612 10260 10744 10266
rect 10612 10254 10692 10260
rect 10692 10202 10744 10208
rect 10796 9994 10824 12310
rect 10888 11898 10916 13126
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11218 10916 11630
rect 10980 11354 11008 15302
rect 11072 15094 11100 15370
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11164 13954 11192 15506
rect 11256 14249 11284 15807
rect 11440 15026 11468 18226
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16969 11560 17002
rect 11518 16960 11574 16969
rect 11518 16895 11574 16904
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11532 16114 11560 16390
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11334 14784 11390 14793
rect 11334 14719 11390 14728
rect 11242 14240 11298 14249
rect 11242 14175 11298 14184
rect 11072 13926 11192 13954
rect 11072 12442 11100 13926
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12436 11112 12442
rect 11164 12434 11192 12582
rect 11164 12406 11284 12434
rect 11060 12378 11112 12384
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11164 11898 11192 12310
rect 11256 12306 11284 12406
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10888 10810 10916 11154
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10538 10916 10746
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10876 10124 10928 10130
rect 10980 10112 11008 11154
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10810 11192 10950
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10928 10084 11008 10112
rect 10876 10066 10928 10072
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10888 9722 10916 10066
rect 11072 9926 11100 10610
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11164 10198 11192 10542
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11256 9722 11284 10066
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8673 10272 8842
rect 10230 8664 10286 8673
rect 10230 8599 10286 8608
rect 10140 8492 10192 8498
rect 10192 8452 10456 8480
rect 10140 8434 10192 8440
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 10152 7886 10180 8026
rect 9312 7880 9364 7886
rect 9588 7880 9640 7886
rect 9312 7822 9364 7828
rect 9586 7848 9588 7857
rect 10140 7880 10192 7886
rect 9640 7848 9642 7857
rect 10140 7822 10192 7828
rect 9586 7783 9642 7792
rect 10428 7546 10456 8452
rect 10612 8362 10640 8978
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 6866 9444 7142
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 5914 9168 6054
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9126 4992 9182 5001
rect 9126 4927 9182 4936
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8758 3360 8814 3369
rect 8758 3295 8814 3304
rect 8772 3126 8800 3295
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8956 2961 8984 3878
rect 8942 2952 8998 2961
rect 8942 2887 8998 2896
rect 9048 2514 9076 4558
rect 9140 2774 9168 4927
rect 9232 4554 9260 6258
rect 9324 6254 9352 6598
rect 9416 6254 9444 6802
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 5137 9352 5170
rect 9310 5128 9366 5137
rect 9310 5063 9366 5072
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9324 4622 9352 4762
rect 9416 4690 9444 6190
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3058 9444 3334
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9140 2746 9260 2774
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 8668 1284 8720 1290
rect 8668 1226 8720 1232
rect 8588 1142 8892 1170
rect 8864 800 8892 1142
rect 9232 800 9260 2746
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9324 1494 9352 2382
rect 9508 1562 9536 7414
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10152 6798 10180 7278
rect 10336 7256 10364 7482
rect 10416 7268 10468 7274
rect 10336 7228 10416 7256
rect 10416 7210 10468 7216
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10612 5778 10640 8298
rect 10704 8090 10732 8366
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10796 7392 10824 8774
rect 11164 8498 11192 8978
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10704 7364 10824 7392
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9600 4060 9628 5578
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4282 9812 4558
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9680 4208 9732 4214
rect 9678 4176 9680 4185
rect 9732 4176 9734 4185
rect 9678 4111 9734 4120
rect 9600 4032 9720 4060
rect 9692 3942 9720 4032
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9968 3126 9996 5170
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4486 10364 4966
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4146 10548 4422
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10060 3194 10088 4014
rect 10152 3942 10180 4082
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10704 3738 10732 7364
rect 10888 7002 10916 8298
rect 11256 7954 11284 8842
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7546 11008 7686
rect 11242 7576 11298 7585
rect 10968 7540 11020 7546
rect 11242 7511 11298 7520
rect 10968 7482 11020 7488
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 5642 10824 6666
rect 11072 5914 11100 6938
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 5914 11192 6666
rect 11256 6254 11284 7511
rect 11348 7342 11376 14719
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 11830 11468 13806
rect 11532 12442 11560 16050
rect 11624 15706 11652 21286
rect 11716 18834 11744 24754
rect 12072 23792 12124 23798
rect 12072 23734 12124 23740
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11900 20602 11928 20810
rect 11992 20641 12020 21558
rect 11978 20632 12034 20641
rect 11888 20596 11940 20602
rect 11978 20567 12034 20576
rect 11888 20538 11940 20544
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11900 19378 11928 19654
rect 12084 19446 12112 23734
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11808 18057 11836 19110
rect 11900 18290 11928 19314
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11992 18057 12020 19110
rect 12176 18986 12204 22918
rect 12268 21486 12296 26726
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12360 22778 12388 26182
rect 12544 25974 12572 29650
rect 12636 29170 12664 30126
rect 12728 29753 12756 30602
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12912 30326 12940 30534
rect 13556 30394 13584 31690
rect 13924 31346 13952 31962
rect 14004 31816 14056 31822
rect 14004 31758 14056 31764
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 13820 30592 13872 30598
rect 13820 30534 13872 30540
rect 13544 30388 13596 30394
rect 13544 30330 13596 30336
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13832 29850 13860 30534
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 12714 29744 12770 29753
rect 12714 29679 12770 29688
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12728 28762 12756 29679
rect 13832 29646 13860 29786
rect 13820 29640 13872 29646
rect 13542 29608 13598 29617
rect 13820 29582 13872 29588
rect 13542 29543 13598 29552
rect 13556 29510 13584 29543
rect 12992 29504 13044 29510
rect 12990 29472 12992 29481
rect 13544 29504 13596 29510
rect 13044 29472 13046 29481
rect 13544 29446 13596 29452
rect 12990 29407 13046 29416
rect 13818 29336 13874 29345
rect 13818 29271 13874 29280
rect 13832 29238 13860 29271
rect 13820 29232 13872 29238
rect 13726 29200 13782 29209
rect 13820 29174 13872 29180
rect 13726 29135 13782 29144
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12716 28756 12768 28762
rect 12716 28698 12768 28704
rect 13452 28484 13504 28490
rect 13452 28426 13504 28432
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 13464 27062 13492 28426
rect 13636 28416 13688 28422
rect 13556 28376 13636 28404
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12636 25226 12664 25978
rect 12808 25764 12860 25770
rect 12808 25706 12860 25712
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 23118 12572 24550
rect 12636 24206 12664 25162
rect 12820 24886 12848 25706
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13372 25378 13400 26794
rect 13452 26512 13504 26518
rect 13452 26454 13504 26460
rect 13280 25350 13400 25378
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 13188 24818 13216 25094
rect 13280 24818 13308 25350
rect 13464 25294 13492 26454
rect 13556 26382 13584 28376
rect 13636 28358 13688 28364
rect 13740 27962 13768 29135
rect 13924 28558 13952 31282
rect 14016 29102 14044 31758
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13648 27934 13768 27962
rect 13648 26602 13676 27934
rect 13728 27872 13780 27878
rect 13728 27814 13780 27820
rect 13740 27606 13768 27814
rect 13728 27600 13780 27606
rect 13728 27542 13780 27548
rect 14016 27402 14044 29038
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13740 26761 13768 27270
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 13726 26752 13782 26761
rect 13726 26687 13782 26696
rect 13648 26574 13768 26602
rect 13636 26512 13688 26518
rect 13636 26454 13688 26460
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13544 26240 13596 26246
rect 13544 26182 13596 26188
rect 13556 25498 13584 26182
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12624 24200 12676 24206
rect 12622 24168 12624 24177
rect 13084 24200 13136 24206
rect 12676 24168 12678 24177
rect 13084 24142 13136 24148
rect 12622 24103 12678 24112
rect 13096 23866 13124 24142
rect 13266 23896 13322 23905
rect 13084 23860 13136 23866
rect 13266 23831 13322 23840
rect 13084 23802 13136 23808
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12636 22094 12664 23462
rect 12820 23322 12848 23598
rect 13280 23594 13308 23831
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 13372 22710 13400 24550
rect 13452 24064 13504 24070
rect 13450 24032 13452 24041
rect 13504 24032 13506 24041
rect 13450 23967 13506 23976
rect 13464 23186 13492 23967
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13556 23066 13584 24822
rect 13464 23038 13584 23066
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13360 22160 13412 22166
rect 13360 22102 13412 22108
rect 12544 22066 12664 22094
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12268 19854 12296 20334
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12084 18958 12204 18986
rect 12084 18630 12112 18958
rect 12268 18698 12296 19654
rect 12360 19242 12388 21354
rect 12438 20224 12494 20233
rect 12438 20159 12494 20168
rect 12452 19990 12480 20159
rect 12544 20058 12572 22066
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 12636 21010 12664 21830
rect 13188 21622 13216 21830
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 13176 21616 13228 21622
rect 13176 21558 13228 21564
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12636 19854 12664 20198
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12544 19334 12572 19790
rect 12452 19306 12572 19334
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12360 18834 12388 19178
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12176 18290 12204 18634
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11794 18048 11850 18057
rect 11794 17983 11850 17992
rect 11978 18048 12034 18057
rect 11978 17983 12034 17992
rect 12084 17542 12112 18158
rect 12360 17882 12388 18566
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11716 17270 11744 17478
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11716 16046 11744 17206
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11900 16969 11928 17002
rect 11886 16960 11942 16969
rect 11886 16895 11942 16904
rect 11992 16590 12020 17138
rect 12084 16726 12112 17478
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11980 16584 12032 16590
rect 11900 16544 11980 16572
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11716 14482 11744 15982
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11808 13938 11836 14758
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11702 13016 11758 13025
rect 11702 12951 11758 12960
rect 11716 12714 11744 12951
rect 11900 12918 11928 16544
rect 11980 16526 12032 16532
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 14482 12020 15846
rect 12084 15570 12112 16662
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12176 15502 12204 17818
rect 12452 17814 12480 19306
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 19122 12756 19178
rect 12544 19094 12756 19122
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12268 16425 12296 16526
rect 12254 16416 12310 16425
rect 12254 16351 12310 16360
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12268 15706 12296 16118
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12164 15496 12216 15502
rect 12084 15444 12164 15450
rect 12084 15438 12216 15444
rect 12084 15422 12204 15438
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11992 14278 12020 14418
rect 12084 14346 12112 15422
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11992 13462 12020 13806
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 13297 12112 13330
rect 12070 13288 12126 13297
rect 12070 13223 12072 13232
rect 12124 13223 12126 13232
rect 12072 13194 12124 13200
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11704 12708 11756 12714
rect 11900 12696 11928 12854
rect 11992 12850 12020 13126
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11900 12668 12020 12696
rect 11704 12650 11756 12656
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11532 11898 11560 12378
rect 11624 12345 11652 12582
rect 11702 12472 11758 12481
rect 11992 12424 12020 12668
rect 11702 12407 11758 12416
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11716 12238 11744 12407
rect 11900 12396 12020 12424
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11426 10432 11482 10441
rect 11532 10418 11560 11698
rect 11624 11286 11652 11766
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11532 10390 11652 10418
rect 11426 10367 11482 10376
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11440 7206 11468 10367
rect 11624 10305 11652 10390
rect 11610 10296 11666 10305
rect 11520 10260 11572 10266
rect 11610 10231 11666 10240
rect 11520 10202 11572 10208
rect 11532 10130 11560 10202
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11532 9382 11560 9862
rect 11624 9450 11652 10066
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11334 6896 11390 6905
rect 11334 6831 11390 6840
rect 11348 6458 11376 6831
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10980 5273 11008 5510
rect 10966 5264 11022 5273
rect 10966 5199 11022 5208
rect 10980 4146 11008 5199
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11058 3768 11114 3777
rect 10692 3732 10744 3738
rect 11058 3703 11114 3712
rect 10692 3674 10744 3680
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9784 1630 9812 2382
rect 9772 1624 9824 1630
rect 9772 1566 9824 1572
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9312 1488 9364 1494
rect 9312 1430 9364 1436
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9600 800 9628 1362
rect 9968 800 9996 2926
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10324 1828 10376 1834
rect 10324 1770 10376 1776
rect 10336 800 10364 1770
rect 10704 800 10732 2858
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10980 1834 11008 2314
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 11072 800 11100 3703
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11440 800 11468 2926
rect 11532 2922 11560 9318
rect 11716 8090 11744 11222
rect 11808 11218 11836 12242
rect 11900 12170 11928 12396
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11900 11898 11928 12106
rect 11992 11937 12020 12242
rect 11978 11928 12034 11937
rect 11888 11892 11940 11898
rect 11978 11863 12034 11872
rect 11888 11834 11940 11840
rect 11900 11354 11928 11834
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11796 10464 11848 10470
rect 11794 10432 11796 10441
rect 11888 10464 11940 10470
rect 11848 10432 11850 10441
rect 11888 10406 11940 10412
rect 11794 10367 11850 10376
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11808 7750 11836 9046
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11624 5234 11652 6326
rect 11808 6254 11836 7142
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11900 5545 11928 10406
rect 11992 7206 12020 11494
rect 12084 10742 12112 13194
rect 12176 12986 12204 15302
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12268 13530 12296 13738
rect 12452 13530 12480 17750
rect 12544 17270 12572 19094
rect 12820 18986 12848 21558
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21078 13400 22102
rect 13464 22098 13492 23038
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13464 20890 13492 22034
rect 13556 22030 13584 22374
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13648 21185 13676 26454
rect 13740 26246 13768 26574
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 13728 26240 13780 26246
rect 13728 26182 13780 26188
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13740 24886 13768 25978
rect 13832 25226 13860 26522
rect 13820 25220 13872 25226
rect 13820 25162 13872 25168
rect 13924 25158 13952 26998
rect 14016 26790 14044 27338
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13728 24880 13780 24886
rect 13728 24822 13780 24828
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13740 22030 13768 24006
rect 13924 23866 13952 24006
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 14004 23792 14056 23798
rect 14002 23760 14004 23769
rect 14056 23760 14058 23769
rect 14002 23695 14058 23704
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13634 21176 13690 21185
rect 13634 21111 13690 21120
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13372 20862 13492 20890
rect 13372 20806 13400 20862
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12912 19378 12940 19994
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 13004 19446 13032 19926
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12728 18958 12848 18986
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 14498 12572 15302
rect 12636 14618 12664 17070
rect 12728 16454 12756 18958
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 13372 18306 13400 20742
rect 13556 19530 13584 21014
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13648 19786 13676 20742
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13556 19502 13676 19530
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13464 18426 13492 19246
rect 13556 18698 13584 19382
rect 13648 18714 13676 19502
rect 13740 19378 13768 20334
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13544 18692 13596 18698
rect 13648 18686 13768 18714
rect 13544 18634 13596 18640
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 12820 17882 12848 18294
rect 13372 18278 13492 18306
rect 13464 18222 13492 18278
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13280 17678 13308 17818
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13372 17592 13400 18158
rect 13452 17604 13504 17610
rect 13372 17564 13452 17592
rect 13452 17546 13504 17552
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15026 12756 15846
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12544 14470 12664 14498
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12176 12481 12204 12650
rect 12162 12472 12218 12481
rect 12162 12407 12218 12416
rect 12268 12238 12296 13330
rect 12360 13025 12388 13330
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12360 12306 12388 12854
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12084 9178 12112 10678
rect 12176 10266 12204 10950
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12268 9722 12296 12038
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12084 8090 12112 8230
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 7886 12204 9658
rect 12360 9042 12388 12038
rect 12452 11098 12480 13262
rect 12544 11898 12572 14282
rect 12636 11898 12664 14470
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12728 11778 12756 14350
rect 12820 13376 12848 17274
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13372 16454 13400 16662
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13096 15978 13124 16390
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15688 13400 16118
rect 13188 15660 13400 15688
rect 13188 15502 13216 15660
rect 13268 15564 13320 15570
rect 13320 15524 13400 15552
rect 13268 15506 13320 15512
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13372 14822 13400 15524
rect 13464 14906 13492 17546
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13556 15026 13584 16118
rect 13648 15570 13676 18566
rect 13740 16096 13768 18686
rect 13832 18358 13860 22034
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13924 18970 13952 19654
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13924 17610 13952 18022
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13924 16794 13952 17138
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14016 16658 14044 19790
rect 14108 17678 14136 41386
rect 14556 38208 14608 38214
rect 14556 38150 14608 38156
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14292 31890 14320 32302
rect 14568 31890 14596 38150
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 14740 32768 14792 32774
rect 14740 32710 14792 32716
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14556 31340 14608 31346
rect 14556 31282 14608 31288
rect 14372 30660 14424 30666
rect 14372 30602 14424 30608
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14200 29714 14228 30126
rect 14188 29708 14240 29714
rect 14188 29650 14240 29656
rect 14384 28150 14412 30602
rect 14568 30394 14596 31282
rect 14556 30388 14608 30394
rect 14556 30330 14608 30336
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14372 28144 14424 28150
rect 14372 28086 14424 28092
rect 14476 27996 14504 28494
rect 14384 27968 14504 27996
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 14200 21350 14228 25162
rect 14292 23497 14320 26726
rect 14278 23488 14334 23497
rect 14278 23423 14334 23432
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14292 22438 14320 23054
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14384 22094 14412 27968
rect 14462 27296 14518 27305
rect 14462 27231 14518 27240
rect 14476 25537 14504 27231
rect 14462 25528 14518 25537
rect 14462 25463 14518 25472
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14476 24342 14504 25298
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14292 22066 14412 22094
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14188 20800 14240 20806
rect 14186 20768 14188 20777
rect 14240 20768 14242 20777
rect 14186 20703 14242 20712
rect 14292 19292 14320 22066
rect 14568 21978 14596 29446
rect 14752 28626 14780 32710
rect 15396 32502 15424 33866
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 15016 32224 15068 32230
rect 15016 32166 15068 32172
rect 15028 31754 15056 32166
rect 15016 31748 15068 31754
rect 15016 31690 15068 31696
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14924 28756 14976 28762
rect 14924 28698 14976 28704
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14660 25430 14688 28154
rect 14936 28014 14964 28698
rect 14924 28008 14976 28014
rect 14924 27950 14976 27956
rect 14740 27328 14792 27334
rect 14738 27296 14740 27305
rect 14832 27328 14884 27334
rect 14792 27296 14794 27305
rect 14832 27270 14884 27276
rect 14738 27231 14794 27240
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14648 25424 14700 25430
rect 14648 25366 14700 25372
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14660 24410 14688 25094
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14646 24032 14702 24041
rect 14646 23967 14702 23976
rect 14660 23730 14688 23967
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14752 22982 14780 25638
rect 14844 25362 14872 27270
rect 15028 26994 15056 29582
rect 15106 29336 15162 29345
rect 15106 29271 15108 29280
rect 15160 29271 15162 29280
rect 15108 29242 15160 29248
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14936 26586 14964 26862
rect 15120 26586 15148 27406
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 15108 26580 15160 26586
rect 15108 26522 15160 26528
rect 15016 26444 15068 26450
rect 15212 26432 15240 30670
rect 15396 30598 15424 32438
rect 15948 31754 15976 42706
rect 16224 33658 16252 53042
rect 16396 50516 16448 50522
rect 16396 50458 16448 50464
rect 16408 41414 16436 50458
rect 16488 50380 16540 50386
rect 16488 50322 16540 50328
rect 16316 41386 16436 41414
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 16224 32842 16252 33594
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 15672 31726 15976 31754
rect 15476 30864 15528 30870
rect 15476 30806 15528 30812
rect 15384 30592 15436 30598
rect 15384 30534 15436 30540
rect 15290 29744 15346 29753
rect 15290 29679 15292 29688
rect 15344 29679 15346 29688
rect 15292 29650 15344 29656
rect 15292 29504 15344 29510
rect 15292 29446 15344 29452
rect 15304 28665 15332 29446
rect 15488 29050 15516 30806
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15580 29306 15608 29990
rect 15568 29300 15620 29306
rect 15568 29242 15620 29248
rect 15396 29022 15516 29050
rect 15290 28656 15346 28665
rect 15290 28591 15346 28600
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15304 27606 15332 28086
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15292 27464 15344 27470
rect 15396 27418 15424 29022
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15488 28490 15516 28902
rect 15476 28484 15528 28490
rect 15476 28426 15528 28432
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15344 27412 15424 27418
rect 15292 27406 15424 27412
rect 15304 27390 15424 27406
rect 15488 26994 15516 27814
rect 15580 26994 15608 29242
rect 15672 29102 15700 31726
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15764 30258 15792 30534
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 15764 30122 15792 30194
rect 15752 30116 15804 30122
rect 15752 30058 15804 30064
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15658 28928 15714 28937
rect 15658 28863 15714 28872
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15016 26386 15068 26392
rect 15120 26404 15240 26432
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14936 25906 14964 26182
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 15028 25226 15056 26386
rect 15120 25906 15148 26404
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 15028 24750 15056 25162
rect 15212 24818 15240 26250
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15396 25702 15424 25978
rect 15476 25832 15528 25838
rect 15476 25774 15528 25780
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 15396 24206 15424 24890
rect 15488 24818 15516 25774
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15384 24200 15436 24206
rect 14830 24168 14886 24177
rect 15384 24142 15436 24148
rect 14830 24103 14886 24112
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14844 22964 14872 24103
rect 15476 23520 15528 23526
rect 15106 23488 15162 23497
rect 15476 23462 15528 23468
rect 15106 23423 15162 23432
rect 15016 23044 15068 23050
rect 14936 23004 15016 23032
rect 14936 22964 14964 23004
rect 15016 22986 15068 22992
rect 14844 22936 14964 22964
rect 14740 22704 14792 22710
rect 14384 21950 14596 21978
rect 14660 22664 14740 22692
rect 14384 20097 14412 21950
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14464 21616 14516 21622
rect 14464 21558 14516 21564
rect 14476 20942 14504 21558
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14370 20088 14426 20097
rect 14370 20023 14426 20032
rect 14476 19922 14504 20878
rect 14568 20874 14596 21830
rect 14660 21622 14688 22664
rect 14844 22692 14872 22936
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 14792 22664 14872 22692
rect 14740 22646 14792 22652
rect 14936 22094 14964 22714
rect 15120 22234 15148 23423
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 14752 22066 14964 22094
rect 15212 22094 15240 23122
rect 15488 22574 15516 23462
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15580 22094 15608 25298
rect 15672 24886 15700 28863
rect 15764 27878 15792 29446
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15752 27396 15804 27402
rect 15752 27338 15804 27344
rect 15764 27062 15792 27338
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15752 26240 15804 26246
rect 15856 26228 15884 30602
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 16026 29472 16082 29481
rect 15948 29238 15976 29446
rect 16026 29407 16082 29416
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15934 28656 15990 28665
rect 16040 28626 16068 29407
rect 16132 29102 16160 29650
rect 16224 29170 16252 31078
rect 16316 30258 16344 41386
rect 16500 33658 16528 50322
rect 16672 41472 16724 41478
rect 16672 41414 16724 41420
rect 16488 33652 16540 33658
rect 16488 33594 16540 33600
rect 16500 32910 16528 33594
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16500 31754 16528 32846
rect 16580 32768 16632 32774
rect 16580 32710 16632 32716
rect 16408 31726 16528 31754
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16316 29646 16344 30194
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16304 29504 16356 29510
rect 16304 29446 16356 29452
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 16120 29096 16172 29102
rect 16120 29038 16172 29044
rect 15934 28591 15936 28600
rect 15988 28591 15990 28600
rect 16028 28620 16080 28626
rect 15936 28562 15988 28568
rect 16028 28562 16080 28568
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 15936 27532 15988 27538
rect 15936 27474 15988 27480
rect 15948 26926 15976 27474
rect 15936 26920 15988 26926
rect 15936 26862 15988 26868
rect 15804 26200 15884 26228
rect 15752 26182 15804 26188
rect 15764 25770 15792 26182
rect 16132 25906 16160 27814
rect 16212 27396 16264 27402
rect 16212 27338 16264 27344
rect 16224 27062 16252 27338
rect 16316 27334 16344 29446
rect 16408 29102 16436 31726
rect 16488 30796 16540 30802
rect 16488 30738 16540 30744
rect 16500 30394 16528 30738
rect 16488 30388 16540 30394
rect 16488 30330 16540 30336
rect 16500 30258 16528 30330
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 16396 29096 16448 29102
rect 16396 29038 16448 29044
rect 16488 29028 16540 29034
rect 16488 28970 16540 28976
rect 16500 27878 16528 28970
rect 16592 28422 16620 32710
rect 16684 32026 16712 41414
rect 16672 32020 16724 32026
rect 16672 31962 16724 31968
rect 16684 30666 16712 31962
rect 16776 31142 16804 53994
rect 17132 53984 17184 53990
rect 17132 53926 17184 53932
rect 17144 45898 17172 53926
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 20364 53106 20392 56200
rect 21744 55214 21772 56200
rect 22374 55448 22430 55457
rect 22374 55383 22430 55392
rect 21744 55186 21864 55214
rect 20352 53100 20404 53106
rect 20352 53042 20404 53048
rect 18972 52964 19024 52970
rect 18972 52906 19024 52912
rect 17224 52488 17276 52494
rect 17224 52430 17276 52436
rect 17132 45892 17184 45898
rect 17132 45834 17184 45840
rect 17236 41414 17264 52430
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 18696 51944 18748 51950
rect 18696 51886 18748 51892
rect 17316 51876 17368 51882
rect 17316 51818 17368 51824
rect 17328 42770 17356 51818
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17316 42764 17368 42770
rect 17316 42706 17368 42712
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 16960 41386 17264 41414
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16776 30734 16804 31078
rect 16764 30728 16816 30734
rect 16764 30670 16816 30676
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16868 30138 16896 32778
rect 16960 31958 16988 41386
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17224 41132 17276 41138
rect 17224 41074 17276 41080
rect 17040 39908 17092 39914
rect 17040 39850 17092 39856
rect 17052 35873 17080 39850
rect 17038 35864 17094 35873
rect 17038 35799 17094 35808
rect 17040 34468 17092 34474
rect 17040 34410 17092 34416
rect 17052 33998 17080 34410
rect 17040 33992 17092 33998
rect 17040 33934 17092 33940
rect 17236 32978 17264 41074
rect 18328 40928 18380 40934
rect 18328 40870 18380 40876
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 18340 38350 18368 40870
rect 18328 38344 18380 38350
rect 18328 38286 18380 38292
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17316 37868 17368 37874
rect 17316 37810 17368 37816
rect 17328 34513 17356 37810
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 18340 34542 18368 34886
rect 18328 34536 18380 34542
rect 17314 34504 17370 34513
rect 18328 34478 18380 34484
rect 17314 34439 17370 34448
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18340 33658 18368 33934
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18420 33516 18472 33522
rect 18420 33458 18472 33464
rect 18432 33114 18460 33458
rect 18420 33108 18472 33114
rect 18420 33050 18472 33056
rect 17224 32972 17276 32978
rect 17224 32914 17276 32920
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 16948 31952 17000 31958
rect 16948 31894 17000 31900
rect 16960 30326 16988 31894
rect 17144 30802 17172 32302
rect 17408 31136 17460 31142
rect 17408 31078 17460 31084
rect 17420 30802 17448 31078
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 17408 30796 17460 30802
rect 17408 30738 17460 30744
rect 16948 30320 17000 30326
rect 16948 30262 17000 30268
rect 16684 30110 16896 30138
rect 16684 28558 16712 30110
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16488 27872 16540 27878
rect 16488 27814 16540 27820
rect 16500 27674 16528 27814
rect 16488 27668 16540 27674
rect 16488 27610 16540 27616
rect 16500 27334 16528 27610
rect 16304 27328 16356 27334
rect 16302 27296 16304 27305
rect 16488 27328 16540 27334
rect 16356 27296 16358 27305
rect 16358 27254 16436 27282
rect 16488 27270 16540 27276
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16302 27231 16358 27240
rect 16212 27056 16264 27062
rect 16212 26998 16264 27004
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 15752 25764 15804 25770
rect 15752 25706 15804 25712
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15672 24410 15700 24822
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15212 22066 15332 22094
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14660 20602 14688 21286
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14660 19922 14688 20538
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14554 19544 14610 19553
rect 14554 19479 14610 19488
rect 14200 19264 14320 19292
rect 14372 19304 14424 19310
rect 14200 19174 14228 19264
rect 14372 19246 14424 19252
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14384 18426 14412 19246
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14188 18080 14240 18086
rect 14186 18048 14188 18057
rect 14240 18048 14242 18057
rect 14186 17983 14242 17992
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14002 16280 14058 16289
rect 14002 16215 14058 16224
rect 14016 16182 14044 16215
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13740 16068 13952 16096
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15570 13768 15846
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13832 15416 13860 15914
rect 13740 15388 13860 15416
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13464 14878 13584 14906
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13188 14074 13216 14554
rect 13372 14074 13400 14758
rect 13464 14278 13492 14758
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13464 13734 13492 13874
rect 13360 13728 13412 13734
rect 13358 13696 13360 13705
rect 13452 13728 13504 13734
rect 13412 13696 13414 13705
rect 13452 13670 13504 13676
rect 12950 13628 13258 13637
rect 13358 13631 13414 13640
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12820 13348 12940 13376
rect 12912 13190 12940 13348
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 12636 11762 12756 11778
rect 13188 11762 13216 12378
rect 13372 11914 13400 13126
rect 13464 12986 13492 13670
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13464 12238 13492 12922
rect 13556 12458 13584 14878
rect 13648 14822 13676 15302
rect 13740 15042 13768 15388
rect 13924 15144 13952 16068
rect 13924 15116 14044 15144
rect 13740 15014 13860 15042
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 13394 13676 14486
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13740 12782 13768 13466
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13740 12617 13768 12718
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13556 12430 13768 12458
rect 13832 12442 13860 15014
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14482 13952 14894
rect 14016 14550 14044 15116
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13636 12368 13688 12374
rect 13634 12336 13636 12345
rect 13688 12336 13690 12345
rect 13740 12322 13768 12430
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13740 12294 13860 12322
rect 13634 12271 13690 12280
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13280 11886 13400 11914
rect 12624 11756 12756 11762
rect 12676 11750 12756 11756
rect 13176 11756 13228 11762
rect 12624 11698 12676 11704
rect 13176 11698 13228 11704
rect 12452 11070 12572 11098
rect 12544 11014 12572 11070
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12636 10792 12664 11698
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11529 12756 11630
rect 13280 11540 13308 11886
rect 13464 11830 13492 12038
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13372 11642 13400 11766
rect 13556 11762 13584 11834
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13372 11614 13584 11642
rect 12714 11520 12770 11529
rect 13280 11512 13492 11540
rect 12714 11455 12770 11464
rect 12728 11286 12756 11455
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13188 11308 13400 11336
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 13084 11280 13136 11286
rect 13188 11268 13216 11308
rect 13136 11240 13216 11268
rect 13084 11222 13136 11228
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12544 10764 12664 10792
rect 12544 10198 12572 10764
rect 13188 10470 13216 11086
rect 13280 10606 13308 11154
rect 13372 11150 13400 11308
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13464 10792 13492 11512
rect 13556 11218 13584 11614
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13648 11393 13676 11562
rect 13634 11384 13690 11393
rect 13634 11319 13690 11328
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13464 10764 13584 10792
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13176 10464 13228 10470
rect 12714 10432 12770 10441
rect 13176 10406 13228 10412
rect 12714 10367 12770 10376
rect 12728 10198 12756 10367
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 13174 9752 13230 9761
rect 13174 9687 13230 9696
rect 12452 9654 12756 9674
rect 12440 9648 12756 9654
rect 12492 9646 12756 9648
rect 12728 9636 12756 9646
rect 12728 9608 12848 9636
rect 12440 9590 12492 9596
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12636 9178 12664 9454
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8673 12296 8842
rect 12254 8664 12310 8673
rect 12452 8634 12480 8910
rect 12254 8599 12310 8608
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11980 6792 12032 6798
rect 12084 6780 12112 7346
rect 12268 6866 12296 7958
rect 12452 7954 12480 8434
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12544 7834 12572 8978
rect 12452 7806 12572 7834
rect 12452 7528 12480 7806
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12360 7500 12480 7528
rect 12360 7410 12388 7500
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12360 7002 12388 7142
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12346 6896 12402 6905
rect 12256 6860 12308 6866
rect 12346 6831 12402 6840
rect 12256 6802 12308 6808
rect 12032 6752 12112 6780
rect 11980 6734 12032 6740
rect 11992 6390 12020 6734
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 11980 6112 12032 6118
rect 12176 6089 12204 6190
rect 11980 6054 12032 6060
rect 12162 6080 12218 6089
rect 11992 5953 12020 6054
rect 12162 6015 12218 6024
rect 11978 5944 12034 5953
rect 11978 5879 12034 5888
rect 11886 5536 11942 5545
rect 11886 5471 11942 5480
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11624 5030 11652 5170
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11794 4584 11850 4593
rect 11794 4519 11850 4528
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11716 2990 11744 3402
rect 11808 3398 11836 4519
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11900 2774 11928 4014
rect 11992 3738 12020 5170
rect 12176 4146 12204 5238
rect 12268 5166 12296 6666
rect 12360 6254 12388 6831
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5953 12388 6054
rect 12346 5944 12402 5953
rect 12346 5879 12402 5888
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12346 4856 12402 4865
rect 12346 4791 12402 4800
rect 12360 4593 12388 4791
rect 12346 4584 12402 4593
rect 12346 4519 12402 4528
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12084 2990 12112 3402
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 11900 2746 12112 2774
rect 11796 2032 11848 2038
rect 11796 1974 11848 1980
rect 12084 1986 12112 2746
rect 12452 2514 12480 7346
rect 12544 6730 12572 7686
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12636 7002 12664 7482
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12622 6896 12678 6905
rect 12622 6831 12624 6840
rect 12676 6831 12678 6840
rect 12624 6802 12676 6808
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12530 6488 12586 6497
rect 12530 6423 12586 6432
rect 12544 6390 12572 6423
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12636 6202 12664 6598
rect 12544 6174 12664 6202
rect 12544 5794 12572 6174
rect 12622 6080 12678 6089
rect 12622 6015 12678 6024
rect 12636 5914 12664 6015
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12544 5766 12664 5794
rect 12636 4049 12664 5766
rect 12728 5166 12756 9318
rect 12820 9110 12848 9608
rect 13188 9518 13216 9687
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 13266 8528 13322 8537
rect 13266 8463 13322 8472
rect 13280 8430 13308 8463
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12820 8129 12848 8298
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12806 8120 12862 8129
rect 12950 8123 13258 8132
rect 12806 8055 12862 8064
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 5846 12848 7686
rect 12912 7274 12940 7890
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13372 6662 13400 10542
rect 13556 10538 13584 10764
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13544 10124 13596 10130
rect 13464 10084 13544 10112
rect 13464 9586 13492 10084
rect 13544 10066 13596 10072
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8362 13492 9318
rect 13556 8362 13584 9930
rect 13648 9178 13676 11018
rect 13740 10044 13768 12106
rect 13832 10606 13860 12294
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13924 10470 13952 14282
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 12170 14044 13806
rect 14108 13530 14136 17614
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 14958 14228 16594
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 15366 14320 16526
rect 14384 16454 14412 17070
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 16046 14412 16390
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 14200 14414 14228 14486
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 14006 14320 14214
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14384 13852 14412 15982
rect 14476 15162 14504 18770
rect 14568 17814 14596 19479
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14752 17134 14780 22066
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15120 21690 15148 21830
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15304 21078 15332 22066
rect 15488 22066 15608 22094
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 15292 21072 15344 21078
rect 15292 21014 15344 21020
rect 14830 20632 14886 20641
rect 14830 20567 14886 20576
rect 14844 18358 14872 20567
rect 14832 18352 14884 18358
rect 14832 18294 14884 18300
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14292 13824 14412 13852
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14108 13258 14136 13466
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14200 12646 14228 12922
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14292 12434 14320 13824
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14108 12406 14320 12434
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13832 10146 13860 10406
rect 13832 10118 13952 10146
rect 13820 10056 13872 10062
rect 13740 10016 13820 10044
rect 13740 9450 13768 10016
rect 13820 9998 13872 10004
rect 13818 9752 13874 9761
rect 13818 9687 13874 9696
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13832 9042 13860 9687
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13648 8566 13676 8774
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13542 8120 13598 8129
rect 13542 8055 13598 8064
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 13372 5710 13400 6054
rect 13464 5794 13492 7890
rect 13556 7750 13584 8055
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13542 6488 13598 6497
rect 13542 6423 13598 6432
rect 13556 6322 13584 6423
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13542 5944 13598 5953
rect 13542 5879 13544 5888
rect 13596 5879 13598 5888
rect 13544 5850 13596 5856
rect 13648 5794 13676 8366
rect 13740 5914 13768 8774
rect 13924 8634 13952 10118
rect 14016 9722 14044 11698
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9042 14044 9386
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13832 8430 13860 8570
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7886 13952 8230
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13832 6254 13860 7754
rect 13924 6730 13952 7822
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 14016 6458 14044 6802
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13464 5766 13584 5794
rect 13648 5766 13768 5794
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5302 13400 5510
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13004 5030 13032 5102
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 12820 4622 12848 4966
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 13464 4146 13492 4966
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 12622 4040 12678 4049
rect 12622 3975 12678 3984
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12636 3738 12664 3878
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12728 3602 12756 3878
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12544 2446 12572 2926
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 11808 800 11836 1974
rect 12084 1958 12204 1986
rect 12176 800 12204 1958
rect 12544 1737 12572 2382
rect 12530 1728 12586 1737
rect 12820 1714 12848 3538
rect 13372 3194 13400 4082
rect 13450 3904 13506 3913
rect 13450 3839 13506 3848
rect 13464 3534 13492 3839
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13372 2650 13400 2994
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 1686 12940 1714
rect 12530 1663 12586 1672
rect 12452 870 12572 898
rect 6184 128 6236 134
rect 6184 70 6236 76
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12452 202 12480 870
rect 12544 800 12572 870
rect 12912 800 12940 1686
rect 13280 800 13308 2314
rect 13556 2009 13584 5766
rect 13740 4486 13768 5766
rect 13924 5574 13952 6394
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13910 4992 13966 5001
rect 13910 4927 13966 4936
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13542 2000 13598 2009
rect 13542 1935 13598 1944
rect 13648 800 13676 2926
rect 13924 1766 13952 4927
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 1760 13964 1766
rect 13912 1702 13964 1708
rect 14016 800 14044 3538
rect 14108 2553 14136 12406
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11694 14228 12038
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14292 11506 14320 11834
rect 14384 11762 14412 12854
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14200 11478 14320 11506
rect 14200 10282 14228 11478
rect 14476 11354 14504 14350
rect 14568 11898 14596 16662
rect 14660 15502 14688 16934
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14660 14550 14688 14894
rect 14752 14822 14780 16934
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 16250 14872 16458
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14830 15192 14886 15201
rect 14830 15127 14886 15136
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14844 14346 14872 15127
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14844 14006 14872 14282
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14660 12646 14688 13806
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14844 12442 14872 12718
rect 14936 12442 14964 21014
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15028 18970 15056 20198
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 19310 15148 19722
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15212 18766 15240 19450
rect 15304 19145 15332 19790
rect 15384 19168 15436 19174
rect 15290 19136 15346 19145
rect 15384 19110 15436 19116
rect 15290 19071 15346 19080
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15016 18624 15068 18630
rect 15396 18612 15424 19110
rect 15016 18566 15068 18572
rect 15106 18592 15162 18601
rect 15028 17202 15056 18566
rect 15106 18527 15162 18536
rect 15212 18584 15424 18612
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15028 15910 15056 16118
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15120 15858 15148 18527
rect 15212 17882 15240 18584
rect 15488 18290 15516 22066
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15304 17882 15332 18226
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15488 17542 15516 18226
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15474 17368 15530 17377
rect 15580 17338 15608 19654
rect 15474 17303 15530 17312
rect 15568 17332 15620 17338
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15212 16182 15240 16458
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15290 16008 15346 16017
rect 15290 15943 15292 15952
rect 15344 15943 15346 15952
rect 15292 15914 15344 15920
rect 15120 15830 15424 15858
rect 15198 15600 15254 15609
rect 15198 15535 15254 15544
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15028 14958 15056 15302
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 15212 14770 15240 15535
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15120 14742 15240 14770
rect 15120 14328 15148 14742
rect 15028 14300 15148 14328
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14924 12436 14976 12442
rect 15028 12434 15056 14300
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15212 13841 15240 14010
rect 15198 13832 15254 13841
rect 15198 13767 15254 13776
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15120 12646 15148 13126
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15028 12406 15148 12434
rect 14924 12378 14976 12384
rect 14660 12170 14688 12378
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14384 11234 14412 11290
rect 14660 11234 14688 11834
rect 14384 11206 14688 11234
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10470 14320 10542
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14200 10266 14320 10282
rect 14200 10260 14332 10266
rect 14200 10254 14280 10260
rect 14280 10202 14332 10208
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14200 9450 14228 10134
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14186 9344 14242 9353
rect 14186 9279 14242 9288
rect 14200 9042 14228 9279
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 14200 7750 14228 8842
rect 14292 7834 14320 10202
rect 14384 10198 14412 10678
rect 14568 10606 14596 11018
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14462 10296 14518 10305
rect 14462 10231 14518 10240
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14384 9353 14412 9522
rect 14370 9344 14426 9353
rect 14370 9279 14426 9288
rect 14476 9058 14504 10231
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14384 9042 14504 9058
rect 14384 9036 14516 9042
rect 14384 9030 14464 9036
rect 14384 8634 14412 9030
rect 14464 8978 14516 8984
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14384 8362 14412 8570
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14476 8129 14504 8298
rect 14462 8120 14518 8129
rect 14462 8055 14518 8064
rect 14292 7806 14504 7834
rect 14188 7744 14240 7750
rect 14280 7744 14332 7750
rect 14188 7686 14240 7692
rect 14278 7712 14280 7721
rect 14332 7712 14334 7721
rect 14278 7647 14334 7656
rect 14476 6848 14504 7806
rect 14384 6820 14504 6848
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 6322 14320 6598
rect 14384 6390 14412 6820
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14384 5846 14412 6326
rect 14568 6322 14596 9862
rect 14660 9654 14688 11206
rect 14752 9994 14780 12174
rect 14936 12073 14964 12378
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15028 12102 15056 12242
rect 15120 12238 15148 12406
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15016 12096 15068 12102
rect 14922 12064 14978 12073
rect 15016 12038 15068 12044
rect 14922 11999 14978 12008
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14844 11336 14872 11698
rect 15028 11626 15056 12038
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15016 11348 15068 11354
rect 14844 11308 15016 11336
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14844 11082 14872 11154
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14936 10470 14964 11308
rect 15016 11290 15068 11296
rect 15120 11200 15148 12174
rect 15028 11172 15148 11200
rect 15028 10742 15056 11172
rect 15212 11098 15240 13126
rect 15304 11218 15332 14962
rect 15396 14090 15424 15830
rect 15488 14278 15516 17303
rect 15568 17274 15620 17280
rect 15566 15600 15622 15609
rect 15566 15535 15622 15544
rect 15580 15502 15608 15535
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15580 15162 15608 15438
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15580 14618 15608 15098
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15396 14062 15516 14090
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15396 13274 15424 13738
rect 15488 13569 15516 14062
rect 15474 13560 15530 13569
rect 15474 13495 15530 13504
rect 15396 13258 15516 13274
rect 15396 13252 15528 13258
rect 15396 13246 15476 13252
rect 15476 13194 15528 13200
rect 15580 13190 15608 14418
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15396 12102 15424 13126
rect 15474 13016 15530 13025
rect 15474 12951 15530 12960
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15120 11070 15240 11098
rect 15292 11076 15344 11082
rect 15120 11014 15148 11070
rect 15292 11018 15344 11024
rect 15108 11008 15160 11014
rect 15304 10962 15332 11018
rect 15108 10950 15160 10956
rect 15212 10934 15332 10962
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14844 9926 14872 10406
rect 14936 10305 14964 10406
rect 14922 10296 14978 10305
rect 14922 10231 14978 10240
rect 15120 10146 15148 10406
rect 14936 10118 15148 10146
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14660 8566 14688 9590
rect 14832 9512 14884 9518
rect 14936 9500 14964 10118
rect 15212 9674 15240 10934
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15120 9646 15240 9674
rect 15120 9518 15148 9646
rect 14884 9472 14964 9500
rect 15108 9512 15160 9518
rect 14832 9454 14884 9460
rect 15108 9454 15160 9460
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14660 7954 14688 8366
rect 14752 8362 14780 9386
rect 14844 8362 14872 9454
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 5234 14504 5510
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14278 4856 14334 4865
rect 14278 4791 14334 4800
rect 14292 4214 14320 4791
rect 14384 4282 14412 5034
rect 14476 4282 14504 5170
rect 14568 4758 14596 6258
rect 14660 5166 14688 7686
rect 14738 6624 14794 6633
rect 14738 6559 14794 6568
rect 14752 5846 14780 6559
rect 14844 6458 14872 8298
rect 14936 7954 14964 8978
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15120 8634 15148 8774
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15212 8430 15240 8774
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15304 8022 15332 10746
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14922 6896 14978 6905
rect 14922 6831 14978 6840
rect 14936 6730 14964 6831
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 15016 6656 15068 6662
rect 14922 6624 14978 6633
rect 15016 6598 15068 6604
rect 14922 6559 14978 6568
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14752 5710 14780 5782
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14738 5536 14794 5545
rect 14738 5471 14794 5480
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14752 4486 14780 5471
rect 14936 5409 14964 6559
rect 15028 6458 15056 6598
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15120 6304 15148 7754
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6798 15240 7142
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15028 6276 15148 6304
rect 14922 5400 14978 5409
rect 14922 5335 14978 5344
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 4690 14872 4966
rect 14936 4758 14964 5034
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14660 4078 14688 4422
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14462 3768 14518 3777
rect 14462 3703 14518 3712
rect 14476 3534 14504 3703
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14094 2544 14150 2553
rect 14094 2479 14150 2488
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 1902 14136 2246
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 14384 800 14412 2450
rect 14752 800 14780 2926
rect 15028 2774 15056 6276
rect 15212 6254 15240 6734
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 6390 15332 6598
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5370 15148 5578
rect 15212 5370 15240 5782
rect 15396 5658 15424 12038
rect 15488 11082 15516 12951
rect 15566 12608 15622 12617
rect 15566 12543 15622 12552
rect 15580 12306 15608 12543
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15488 8362 15516 10610
rect 15580 9042 15608 11834
rect 15672 10690 15700 24346
rect 15764 19242 15792 25706
rect 16118 25392 16174 25401
rect 16118 25327 16174 25336
rect 16132 25294 16160 25327
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 16040 23866 16068 25094
rect 16132 24954 16160 25230
rect 16408 25158 16436 27254
rect 16500 27062 16528 27270
rect 16488 27056 16540 27062
rect 16488 26998 16540 27004
rect 16592 26874 16620 27270
rect 16500 26846 16620 26874
rect 16500 25702 16528 26846
rect 16684 26042 16712 28358
rect 16776 27470 16804 29990
rect 16960 29714 16988 30262
rect 17040 30184 17092 30190
rect 17040 30126 17092 30132
rect 16856 29708 16908 29714
rect 16856 29650 16908 29656
rect 16948 29708 17000 29714
rect 16948 29650 17000 29656
rect 16868 29306 16896 29650
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16868 28218 16896 28562
rect 16948 28484 17000 28490
rect 16948 28426 17000 28432
rect 16960 28218 16988 28426
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16868 27538 16896 28154
rect 17052 28082 17080 30126
rect 17224 30116 17276 30122
rect 17224 30058 17276 30064
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16868 26994 16896 27474
rect 17144 26994 17172 29582
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16776 26382 16804 26726
rect 17130 26480 17186 26489
rect 17130 26415 17186 26424
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16408 24970 16436 25094
rect 16408 24954 16528 24970
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 16304 24948 16356 24954
rect 16408 24948 16540 24954
rect 16408 24942 16488 24948
rect 16304 24890 16356 24896
rect 16488 24890 16540 24896
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22710 15884 22918
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15750 17912 15806 17921
rect 15750 17847 15752 17856
rect 15804 17847 15806 17856
rect 15752 17818 15804 17824
rect 15764 17678 15792 17818
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15856 16046 15884 20198
rect 15948 17746 15976 23122
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16132 22098 16160 22918
rect 16224 22778 16252 24754
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16132 21554 16160 22034
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16316 21434 16344 24890
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16500 24614 16528 24686
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16500 23769 16528 24550
rect 16486 23760 16542 23769
rect 16486 23695 16542 23704
rect 16394 23624 16450 23633
rect 16394 23559 16450 23568
rect 16408 22681 16436 23559
rect 16500 23254 16528 23695
rect 16488 23248 16540 23254
rect 16488 23190 16540 23196
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16394 22672 16450 22681
rect 16394 22607 16450 22616
rect 16396 22568 16448 22574
rect 16394 22536 16396 22545
rect 16448 22536 16450 22545
rect 16394 22471 16450 22480
rect 16224 21406 16344 21434
rect 16394 21448 16450 21457
rect 16224 19446 16252 21406
rect 16394 21383 16450 21392
rect 16408 21350 16436 21383
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16316 21010 16344 21286
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16316 20262 16344 20810
rect 16408 20398 16436 21014
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18154 16068 18566
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15948 17490 15976 17682
rect 15948 17462 16068 17490
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15764 14550 15792 15982
rect 15948 15978 15976 17274
rect 16040 16726 16068 17462
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 16118 16688 16174 16697
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15948 15337 15976 15370
rect 16040 15366 16068 16662
rect 16118 16623 16174 16632
rect 16028 15360 16080 15366
rect 15934 15328 15990 15337
rect 16028 15302 16080 15308
rect 15934 15263 15990 15272
rect 16132 14890 16160 16623
rect 16224 16250 16252 19110
rect 16316 18057 16344 19110
rect 16408 18902 16436 19314
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 16500 18834 16528 22918
rect 16592 22030 16620 25638
rect 16684 24070 16712 25774
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 22982 16712 24006
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16684 21690 16712 22578
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16776 21026 16804 25162
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16868 22778 16896 23666
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16868 21554 16896 22442
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16684 20998 16804 21026
rect 16684 20058 16712 20998
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 20058 16804 20878
rect 16868 20466 16896 21490
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16868 18290 16896 20402
rect 16960 19786 16988 24550
rect 17144 24342 17172 26415
rect 17132 24336 17184 24342
rect 17132 24278 17184 24284
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17052 20942 17080 24210
rect 17236 24070 17264 30058
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 17408 29572 17460 29578
rect 17408 29514 17460 29520
rect 17328 28626 17356 29514
rect 17420 29238 17448 29514
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 17512 28937 17540 29990
rect 17498 28928 17554 28937
rect 17498 28863 17554 28872
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17328 24750 17356 28358
rect 17604 27470 17632 32846
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18432 32502 18460 32710
rect 18420 32496 18472 32502
rect 18420 32438 18472 32444
rect 18432 31754 18460 32438
rect 18524 32366 18552 33798
rect 18708 33114 18736 51886
rect 18788 49428 18840 49434
rect 18788 49370 18840 49376
rect 18800 41414 18828 49370
rect 18800 41386 18920 41414
rect 18696 33108 18748 33114
rect 18616 33068 18696 33096
rect 18616 32842 18644 33068
rect 18696 33050 18748 33056
rect 18788 32904 18840 32910
rect 18788 32846 18840 32852
rect 18604 32836 18656 32842
rect 18604 32778 18656 32784
rect 18512 32360 18564 32366
rect 18512 32302 18564 32308
rect 18432 31726 18552 31754
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17880 30326 17908 31282
rect 18420 30592 18472 30598
rect 18420 30534 18472 30540
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 17868 30320 17920 30326
rect 17868 30262 17920 30268
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18340 29510 18368 30126
rect 18432 29578 18460 30534
rect 18524 29866 18552 31726
rect 18616 30841 18644 32778
rect 18800 31958 18828 32846
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 18696 31748 18748 31754
rect 18696 31690 18748 31696
rect 18602 30832 18658 30841
rect 18602 30767 18658 30776
rect 18708 30666 18736 31690
rect 18696 30660 18748 30666
rect 18696 30602 18748 30608
rect 18524 29838 18644 29866
rect 18512 29776 18564 29782
rect 18512 29718 18564 29724
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18340 29152 18368 29446
rect 18248 29124 18368 29152
rect 18248 29034 18276 29124
rect 17960 29028 18012 29034
rect 17960 28970 18012 28976
rect 18236 29028 18288 29034
rect 18236 28970 18288 28976
rect 18328 29028 18380 29034
rect 18328 28970 18380 28976
rect 17776 28960 17828 28966
rect 17776 28902 17828 28908
rect 17788 28558 17816 28902
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 17144 21457 17172 21558
rect 17130 21448 17186 21457
rect 17130 21383 17186 21392
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 17038 19408 17094 19417
rect 17038 19343 17094 19352
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16302 18048 16358 18057
rect 16302 17983 16358 17992
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 16408 17513 16436 17546
rect 16764 17536 16816 17542
rect 16394 17504 16450 17513
rect 16764 17478 16816 17484
rect 16394 17439 16450 17448
rect 16408 16697 16436 17439
rect 16394 16688 16450 16697
rect 16304 16652 16356 16658
rect 16394 16623 16450 16632
rect 16304 16594 16356 16600
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16224 15706 16252 15914
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16316 15570 16344 16594
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16408 15162 16436 16050
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15856 13682 15884 14826
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 13802 15976 14350
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16040 13870 16068 14282
rect 16224 14278 16252 14894
rect 16500 14328 16528 16186
rect 16684 16153 16712 16390
rect 16670 16144 16726 16153
rect 16670 16079 16726 16088
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16592 14618 16620 14962
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16316 14300 16528 14328
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 16224 13734 16252 14214
rect 15764 13654 15884 13682
rect 16028 13728 16080 13734
rect 16212 13728 16264 13734
rect 16028 13670 16080 13676
rect 16118 13696 16174 13705
rect 15764 10810 15792 13654
rect 15842 13560 15898 13569
rect 16040 13530 16068 13670
rect 16212 13670 16264 13676
rect 16118 13631 16174 13640
rect 15842 13495 15898 13504
rect 16028 13524 16080 13530
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15672 10662 15792 10690
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15580 8566 15608 8978
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15476 6656 15528 6662
rect 15474 6624 15476 6633
rect 15528 6624 15530 6633
rect 15474 6559 15530 6568
rect 15474 6488 15530 6497
rect 15474 6423 15530 6432
rect 15488 6390 15516 6423
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15580 6254 15608 7414
rect 15672 7410 15700 9862
rect 15764 8650 15792 10662
rect 15856 10266 15884 13495
rect 16028 13466 16080 13472
rect 16132 13394 16160 13631
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15856 9654 15884 10202
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15948 9178 15976 13262
rect 16040 11898 16068 13330
rect 16118 13016 16174 13025
rect 16118 12951 16174 12960
rect 16132 12782 16160 12951
rect 16224 12850 16252 13670
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16316 11778 16344 14300
rect 16394 14240 16450 14249
rect 16394 14175 16450 14184
rect 16408 13938 16436 14175
rect 16486 14104 16542 14113
rect 16486 14039 16542 14048
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16408 12481 16436 13874
rect 16500 13841 16528 14039
rect 16486 13832 16542 13841
rect 16486 13767 16542 13776
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16592 12986 16620 13670
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16394 12472 16450 12481
rect 16394 12407 16450 12416
rect 16486 12200 16542 12209
rect 16486 12135 16542 12144
rect 16028 11756 16080 11762
rect 16316 11750 16436 11778
rect 16028 11698 16080 11704
rect 16040 11286 16068 11698
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16040 10606 16068 10746
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16040 9353 16068 10542
rect 16132 9926 16160 11222
rect 16224 11218 16252 11494
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16316 11150 16344 11494
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16302 10976 16358 10985
rect 16302 10911 16358 10920
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16224 9738 16252 10678
rect 16132 9710 16252 9738
rect 16316 9738 16344 10911
rect 16408 10674 16436 11750
rect 16500 10742 16528 12135
rect 16592 12073 16620 12582
rect 16578 12064 16634 12073
rect 16578 11999 16634 12008
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16408 9897 16436 9930
rect 16394 9888 16450 9897
rect 16394 9823 16450 9832
rect 16316 9710 16436 9738
rect 16132 9450 16160 9710
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16026 9344 16082 9353
rect 16026 9279 16082 9288
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 15764 8622 15884 8650
rect 15750 8528 15806 8537
rect 15750 8463 15806 8472
rect 15764 8430 15792 8463
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5817 15608 6054
rect 15566 5808 15622 5817
rect 15566 5743 15622 5752
rect 15396 5630 15608 5658
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15304 5030 15332 5170
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 15120 3369 15148 3402
rect 15106 3360 15162 3369
rect 15106 3295 15162 3304
rect 14936 2746 15056 2774
rect 14936 2310 14964 2746
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 15120 800 15148 2450
rect 15304 1465 15332 4966
rect 15488 4826 15516 4966
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15290 1456 15346 1465
rect 15290 1391 15346 1400
rect 15488 800 15516 3538
rect 15580 2378 15608 5630
rect 15672 4214 15700 6666
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15764 3942 15792 6802
rect 15856 6633 15884 8622
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15948 8401 15976 8434
rect 15934 8392 15990 8401
rect 15934 8327 15990 8336
rect 15948 7410 15976 8327
rect 15936 7404 15988 7410
rect 16040 7392 16068 9046
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16132 7460 16160 8910
rect 16224 8838 16252 9590
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16224 8430 16252 8502
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16224 7954 16252 8366
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16212 7472 16264 7478
rect 16132 7432 16212 7460
rect 16212 7414 16264 7420
rect 16040 7364 16160 7392
rect 15936 7346 15988 7352
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 15934 6896 15990 6905
rect 15934 6831 15936 6840
rect 15988 6831 15990 6840
rect 15936 6802 15988 6808
rect 15842 6624 15898 6633
rect 15842 6559 15898 6568
rect 15842 6488 15898 6497
rect 15842 6423 15898 6432
rect 15856 6254 15884 6423
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15856 4282 15884 6190
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5370 15976 6122
rect 16040 5710 16068 7210
rect 16132 6730 16160 7364
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3534 15792 3878
rect 15948 3738 15976 4762
rect 16040 4690 16068 5646
rect 16132 4690 16160 6190
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16040 3942 16068 4218
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15856 800 15884 2926
rect 15948 2378 15976 3674
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 16040 2310 16068 3878
rect 16132 2922 16160 4626
rect 16224 3534 16252 7142
rect 16316 5234 16344 9386
rect 16408 8888 16436 9710
rect 16500 9042 16528 10474
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16488 8900 16540 8906
rect 16408 8860 16488 8888
rect 16488 8842 16540 8848
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7206 16436 7890
rect 16592 7750 16620 11183
rect 16684 8838 16712 14418
rect 16776 11150 16804 17478
rect 16868 16658 16896 18226
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16960 16998 16988 17478
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16854 16144 16910 16153
rect 16854 16079 16910 16088
rect 16868 15910 16896 16079
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 14414 16896 15302
rect 16856 14408 16908 14414
rect 17052 14362 17080 19343
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 18358 17172 18566
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 16454 17172 17478
rect 17236 16794 17264 24006
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17328 17542 17356 20742
rect 17420 19334 17448 26998
rect 17604 26042 17632 27406
rect 17592 26036 17644 26042
rect 17592 25978 17644 25984
rect 17604 25378 17632 25978
rect 17604 25350 17724 25378
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 17512 24206 17540 24890
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17512 22030 17540 22510
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 20641 17540 21966
rect 17498 20632 17554 20641
rect 17604 20602 17632 25230
rect 17696 24954 17724 25350
rect 17684 24948 17736 24954
rect 17684 24890 17736 24896
rect 17788 22094 17816 28494
rect 17972 28404 18000 28970
rect 17880 28376 18000 28404
rect 17880 28150 17908 28376
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17868 28144 17920 28150
rect 17868 28086 17920 28092
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17880 26450 17908 26930
rect 18340 26518 18368 28970
rect 18432 28150 18460 29514
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 18328 26512 18380 26518
rect 18328 26454 18380 26460
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 18420 26308 18472 26314
rect 18420 26250 18472 26256
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18432 26042 18460 26250
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18050 25800 18106 25809
rect 18050 25735 18052 25744
rect 18104 25735 18106 25744
rect 18052 25706 18104 25712
rect 18524 25226 18552 29718
rect 18616 28490 18644 29838
rect 18694 29608 18750 29617
rect 18694 29543 18750 29552
rect 18708 29170 18736 29543
rect 18696 29164 18748 29170
rect 18696 29106 18748 29112
rect 18696 29028 18748 29034
rect 18696 28970 18748 28976
rect 18604 28484 18656 28490
rect 18604 28426 18656 28432
rect 18616 27674 18644 28426
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18616 26246 18644 27406
rect 18708 26489 18736 28970
rect 18800 28626 18828 31894
rect 18892 31754 18920 41386
rect 18984 33114 19012 52906
rect 20444 46980 20496 46986
rect 20444 46922 20496 46928
rect 20812 46980 20864 46986
rect 20812 46922 20864 46928
rect 19708 46436 19760 46442
rect 19708 46378 19760 46384
rect 19064 44192 19116 44198
rect 19064 44134 19116 44140
rect 19076 34626 19104 44134
rect 19432 43784 19484 43790
rect 19432 43726 19484 43732
rect 19156 35692 19208 35698
rect 19156 35634 19208 35640
rect 19168 34746 19196 35634
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 19076 34598 19196 34626
rect 18972 33108 19024 33114
rect 18972 33050 19024 33056
rect 18892 31726 19012 31754
rect 18984 30258 19012 31726
rect 19064 30320 19116 30326
rect 19064 30262 19116 30268
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18892 29510 18920 30194
rect 18972 30116 19024 30122
rect 18972 30058 19024 30064
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18788 28620 18840 28626
rect 18788 28562 18840 28568
rect 18786 27568 18842 27577
rect 18786 27503 18842 27512
rect 18800 27334 18828 27503
rect 18788 27328 18840 27334
rect 18788 27270 18840 27276
rect 18694 26480 18750 26489
rect 18694 26415 18750 26424
rect 18800 26382 18828 27270
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18708 25498 18736 26318
rect 18788 25900 18840 25906
rect 18788 25842 18840 25848
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18340 24750 18368 25094
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18510 24712 18566 24721
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17696 22066 17816 22094
rect 17696 20806 17724 22066
rect 17880 21962 17908 22918
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18340 22710 18368 24686
rect 18420 24676 18472 24682
rect 18510 24647 18512 24656
rect 18420 24618 18472 24624
rect 18564 24647 18566 24656
rect 18512 24618 18564 24624
rect 18432 24206 18460 24618
rect 18420 24200 18472 24206
rect 18616 24154 18644 24890
rect 18696 24880 18748 24886
rect 18696 24822 18748 24828
rect 18420 24142 18472 24148
rect 18524 24126 18644 24154
rect 18524 24070 18552 24126
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 18248 22094 18276 22646
rect 18432 22094 18460 24006
rect 18524 23866 18552 24006
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18248 22066 18368 22094
rect 18432 22066 18552 22094
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17682 20632 17738 20641
rect 17498 20567 17554 20576
rect 17592 20596 17644 20602
rect 17682 20567 17738 20576
rect 17592 20538 17644 20544
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17512 20058 17540 20470
rect 17696 20262 17724 20567
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17590 19816 17646 19825
rect 17512 19514 17540 19790
rect 17590 19751 17646 19760
rect 17604 19718 17632 19751
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17420 19306 17540 19334
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17512 17134 17540 19306
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17500 17128 17552 17134
rect 17328 17076 17500 17082
rect 17328 17070 17552 17076
rect 17328 17054 17540 17070
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17236 16590 17264 16730
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 16856 14350 16908 14356
rect 16868 14249 16896 14350
rect 16960 14334 17080 14362
rect 16854 14240 16910 14249
rect 16854 14175 16910 14184
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16776 10062 16804 10610
rect 16868 10198 16896 13126
rect 16960 12238 16988 14334
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9926 16804 9998
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16948 9648 17000 9654
rect 16946 9616 16948 9625
rect 17000 9616 17002 9625
rect 16946 9551 17002 9560
rect 17052 9466 17080 13398
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17144 10266 17172 12718
rect 17236 12442 17264 12718
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17328 12102 17356 17054
rect 17512 16998 17540 17054
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17222 11792 17278 11801
rect 17222 11727 17278 11736
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17236 9722 17264 11727
rect 17328 10606 17356 12038
rect 17420 11898 17448 16934
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17512 14346 17540 16623
rect 17604 15366 17632 17682
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17696 14958 17724 20198
rect 17788 18766 17816 21830
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18340 20754 18368 22066
rect 18340 20726 18460 20754
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18326 20088 18382 20097
rect 18236 20052 18288 20058
rect 18326 20023 18328 20032
rect 18236 19994 18288 20000
rect 18380 20023 18382 20032
rect 18328 19994 18380 20000
rect 18248 19700 18276 19994
rect 18248 19672 18368 19700
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18340 19394 18368 19672
rect 18248 19366 18368 19394
rect 18432 19378 18460 20726
rect 18524 19854 18552 22066
rect 18616 21690 18644 23122
rect 18708 22778 18736 24822
rect 18800 24070 18828 25842
rect 18892 25838 18920 29446
rect 18984 26790 19012 30058
rect 19076 29209 19104 30262
rect 19168 30054 19196 34598
rect 19444 34066 19472 43726
rect 19720 41414 19748 46378
rect 20168 45892 20220 45898
rect 20168 45834 20220 45840
rect 19720 41386 19840 41414
rect 19524 35080 19576 35086
rect 19524 35022 19576 35028
rect 19432 34060 19484 34066
rect 19432 34002 19484 34008
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 19260 31754 19288 33254
rect 19352 33114 19380 33458
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19444 32910 19472 33390
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19444 32366 19472 32846
rect 19432 32360 19484 32366
rect 19432 32302 19484 32308
rect 19444 32026 19472 32302
rect 19536 32230 19564 35022
rect 19616 34944 19668 34950
rect 19616 34886 19668 34892
rect 19628 34610 19656 34886
rect 19708 34740 19760 34746
rect 19708 34682 19760 34688
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 19524 32224 19576 32230
rect 19524 32166 19576 32172
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19444 31822 19472 31962
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19720 31754 19748 34682
rect 19260 31726 19380 31754
rect 19352 31362 19380 31726
rect 19708 31748 19760 31754
rect 19708 31690 19760 31696
rect 19812 31634 19840 41386
rect 20076 38480 20128 38486
rect 20076 38422 20128 38428
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19892 34400 19944 34406
rect 19892 34342 19944 34348
rect 19720 31606 19840 31634
rect 19720 31482 19748 31606
rect 19708 31476 19760 31482
rect 19708 31418 19760 31424
rect 19352 31334 19840 31362
rect 19616 31272 19668 31278
rect 19616 31214 19668 31220
rect 19708 31272 19760 31278
rect 19708 31214 19760 31220
rect 19524 31136 19576 31142
rect 19524 31078 19576 31084
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19168 29832 19196 29990
rect 19168 29804 19288 29832
rect 19156 29708 19208 29714
rect 19156 29650 19208 29656
rect 19062 29200 19118 29209
rect 19062 29135 19118 29144
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 19064 26784 19116 26790
rect 19064 26726 19116 26732
rect 18972 26376 19024 26382
rect 18970 26344 18972 26353
rect 19024 26344 19026 26353
rect 18970 26279 19026 26288
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 19076 25294 19104 26726
rect 19168 25498 19196 29650
rect 19260 28966 19288 29804
rect 19352 29782 19380 29990
rect 19340 29776 19392 29782
rect 19340 29718 19392 29724
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19352 28218 19380 29514
rect 19536 28558 19564 31078
rect 19628 30258 19656 31214
rect 19720 30734 19748 31214
rect 19708 30728 19760 30734
rect 19708 30670 19760 30676
rect 19812 30546 19840 31334
rect 19720 30518 19840 30546
rect 19616 30252 19668 30258
rect 19616 30194 19668 30200
rect 19616 29504 19668 29510
rect 19616 29446 19668 29452
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19260 27538 19288 27882
rect 19248 27532 19300 27538
rect 19248 27474 19300 27480
rect 19352 27130 19380 28154
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19340 26852 19392 26858
rect 19340 26794 19392 26800
rect 19352 26586 19380 26794
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19524 25900 19576 25906
rect 19524 25842 19576 25848
rect 19536 25498 19564 25842
rect 19156 25492 19208 25498
rect 19156 25434 19208 25440
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19064 25288 19116 25294
rect 19064 25230 19116 25236
rect 19076 24750 19104 25230
rect 19168 24954 19196 25434
rect 19156 24948 19208 24954
rect 19156 24890 19208 24896
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18800 22545 18828 22918
rect 18786 22536 18842 22545
rect 18786 22471 18842 22480
rect 18696 22432 18748 22438
rect 18892 22420 18920 24210
rect 19352 24154 19380 24754
rect 19076 24126 19380 24154
rect 19076 23730 19104 24126
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 19168 23610 19196 24006
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19260 23746 19288 23802
rect 19260 23718 19380 23746
rect 19168 23582 19288 23610
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 18696 22374 18748 22380
rect 18800 22392 18920 22420
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18616 21078 18644 21422
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18420 19372 18472 19378
rect 18248 19242 18276 19366
rect 18420 19314 18472 19320
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18156 18902 18184 19178
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 18156 18612 18184 18838
rect 18248 18680 18276 19178
rect 18340 18902 18368 19246
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18248 18652 18460 18680
rect 18156 18584 18368 18612
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18340 17678 18368 18584
rect 18432 18358 18460 18652
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 18328 17672 18380 17678
rect 18380 17620 18460 17626
rect 18328 17614 18460 17620
rect 17788 17202 17816 17614
rect 18340 17598 18460 17614
rect 17960 17536 18012 17542
rect 17880 17496 17960 17524
rect 17880 17241 17908 17496
rect 17960 17478 18012 17484
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17866 17232 17922 17241
rect 17776 17196 17828 17202
rect 17866 17167 17922 17176
rect 17776 17138 17828 17144
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16232 17908 17070
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17788 16204 17908 16232
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17788 14482 17816 16204
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18248 15434 18276 16118
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18340 15162 18368 17478
rect 18432 17066 18460 17598
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 16114 18460 16594
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18524 16017 18552 19654
rect 18616 18358 18644 20742
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17746 18644 18022
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18510 16008 18566 16017
rect 18420 15972 18472 15978
rect 18510 15943 18566 15952
rect 18420 15914 18472 15920
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18432 15042 18460 15914
rect 18510 15464 18566 15473
rect 18510 15399 18566 15408
rect 18340 15014 18460 15042
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 18248 14414 18276 14758
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17512 12345 17540 14010
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17498 12336 17554 12345
rect 17498 12271 17554 12280
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17512 11354 17540 11834
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17604 10674 17632 13738
rect 17696 13326 17724 14214
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17774 13696 17830 13705
rect 17774 13631 17830 13640
rect 17788 13326 17816 13631
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17880 13190 17908 13874
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17880 12918 17908 13126
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 18156 12714 18184 12922
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18340 12481 18368 15014
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13938 18460 14214
rect 18524 14074 18552 15399
rect 18616 15026 18644 17682
rect 18708 17678 18736 22374
rect 18800 22030 18828 22392
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18800 19922 18828 21286
rect 18892 20806 18920 21830
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18984 21078 19012 21490
rect 19076 21486 19104 22646
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 19168 20874 19196 22714
rect 19260 22234 19288 23582
rect 19352 23186 19380 23718
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19248 22228 19300 22234
rect 19248 22170 19300 22176
rect 19352 22098 19380 23122
rect 19444 22778 19472 24006
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19536 23497 19564 23802
rect 19628 23746 19656 29446
rect 19720 27538 19748 30518
rect 19800 30184 19852 30190
rect 19800 30126 19852 30132
rect 19812 29646 19840 30126
rect 19800 29640 19852 29646
rect 19800 29582 19852 29588
rect 19904 28966 19932 34342
rect 19996 33658 20024 36110
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 19892 28960 19944 28966
rect 19892 28902 19944 28908
rect 20088 28098 20116 38422
rect 20180 35154 20208 45834
rect 20456 36922 20484 46922
rect 20824 43858 20852 46922
rect 21732 46504 21784 46510
rect 21732 46446 21784 46452
rect 20812 43852 20864 43858
rect 20812 43794 20864 43800
rect 21272 43852 21324 43858
rect 21272 43794 21324 43800
rect 21284 43722 21312 43794
rect 21088 43716 21140 43722
rect 21088 43658 21140 43664
rect 21272 43716 21324 43722
rect 21272 43658 21324 43664
rect 20628 43648 20680 43654
rect 21100 43602 21128 43658
rect 20628 43590 20680 43596
rect 20640 41138 20668 43590
rect 21008 43574 21128 43602
rect 21008 41414 21036 43574
rect 21008 41386 21312 41414
rect 20628 41132 20680 41138
rect 20628 41074 20680 41080
rect 21088 38752 21140 38758
rect 21088 38694 21140 38700
rect 20444 36916 20496 36922
rect 20444 36858 20496 36864
rect 20456 35834 20484 36858
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20812 35556 20864 35562
rect 20812 35498 20864 35504
rect 20260 35488 20312 35494
rect 20260 35430 20312 35436
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20168 35148 20220 35154
rect 20168 35090 20220 35096
rect 20180 31754 20208 35090
rect 20272 35086 20300 35430
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20364 32978 20392 34886
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20352 32972 20404 32978
rect 20352 32914 20404 32920
rect 20180 31726 20300 31754
rect 20272 31482 20300 31726
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 20260 31476 20312 31482
rect 20260 31418 20312 31424
rect 20180 30818 20208 31418
rect 20272 30938 20300 31418
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20180 30790 20392 30818
rect 20364 30598 20392 30790
rect 20352 30592 20404 30598
rect 20352 30534 20404 30540
rect 20168 30320 20220 30326
rect 20168 30262 20220 30268
rect 20180 30054 20208 30262
rect 20168 30048 20220 30054
rect 20168 29990 20220 29996
rect 20364 29782 20392 30534
rect 20456 30190 20484 33594
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20536 31680 20588 31686
rect 20536 31622 20588 31628
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20352 29776 20404 29782
rect 20352 29718 20404 29724
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 19812 28070 20116 28098
rect 19708 27532 19760 27538
rect 19708 27474 19760 27480
rect 19708 26444 19760 26450
rect 19708 26386 19760 26392
rect 19720 24818 19748 26386
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19708 24336 19760 24342
rect 19708 24278 19760 24284
rect 19720 23866 19748 24278
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19628 23718 19748 23746
rect 19522 23488 19578 23497
rect 19522 23423 19578 23432
rect 19616 23180 19668 23186
rect 19616 23122 19668 23128
rect 19628 22982 19656 23122
rect 19616 22976 19668 22982
rect 19616 22918 19668 22924
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18970 20496 19026 20505
rect 18970 20431 19026 20440
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18800 17921 18828 18838
rect 18892 18698 18920 19994
rect 18984 19990 19012 20431
rect 18972 19984 19024 19990
rect 19076 19972 19104 20810
rect 19168 20602 19196 20810
rect 19260 20806 19288 21898
rect 19338 21856 19394 21865
rect 19338 21791 19394 21800
rect 19352 21049 19380 21791
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19338 21040 19394 21049
rect 19338 20975 19394 20984
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19352 20602 19380 20975
rect 19444 20913 19472 21286
rect 19430 20904 19486 20913
rect 19430 20839 19486 20848
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19352 20398 19380 20538
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19156 19984 19208 19990
rect 19076 19944 19156 19972
rect 18972 19926 19024 19932
rect 19156 19926 19208 19932
rect 19156 19780 19208 19786
rect 19156 19722 19208 19728
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 19076 19378 19104 19654
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18786 17912 18842 17921
rect 18786 17847 18842 17856
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18708 16561 18736 16594
rect 18694 16552 18750 16561
rect 18892 16522 18920 18226
rect 18694 16487 18750 16496
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18892 16402 18920 16458
rect 18800 16374 18920 16402
rect 18800 16182 18828 16374
rect 18984 16266 19012 19246
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18290 19104 19110
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19062 17776 19118 17785
rect 19062 17711 19064 17720
rect 19116 17711 19118 17720
rect 19064 17682 19116 17688
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18892 16238 19012 16266
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18524 13462 18552 14010
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18326 12472 18382 12481
rect 17684 12436 17736 12442
rect 18326 12407 18382 12416
rect 17684 12378 17736 12384
rect 17696 12073 17724 12378
rect 18432 12186 18460 12922
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18340 12158 18460 12186
rect 17776 12096 17828 12102
rect 17682 12064 17738 12073
rect 17776 12038 17828 12044
rect 17682 11999 17738 12008
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17696 11082 17724 11290
rect 17788 11150 17816 12038
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11778 18368 12158
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18248 11750 18368 11778
rect 17866 11384 17922 11393
rect 17866 11319 17868 11328
rect 17920 11319 17922 11328
rect 17868 11290 17920 11296
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 18248 10996 18276 11750
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 17880 10968 18276 10996
rect 17880 10810 17908 10968
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10062 17724 10406
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17880 10169 17908 10202
rect 17866 10160 17922 10169
rect 17866 10095 17922 10104
rect 18340 10062 18368 11630
rect 18432 10674 18460 12038
rect 18524 11694 18552 12582
rect 18616 11762 18644 12582
rect 18708 12442 18736 15982
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18708 11218 18736 12242
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17224 9716 17276 9722
rect 17880 9704 17908 9862
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17880 9676 18000 9704
rect 17224 9658 17276 9664
rect 17592 9512 17644 9518
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16868 9438 17080 9466
rect 17236 9472 17592 9500
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 8362 16712 8774
rect 16776 8634 16804 9386
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16776 8022 16804 8570
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16486 7576 16542 7585
rect 16486 7511 16542 7520
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16500 6905 16528 7511
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16486 6896 16542 6905
rect 16486 6831 16542 6840
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16408 4146 16436 6258
rect 16500 5370 16528 6326
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16500 4622 16528 4694
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16224 800 16252 2858
rect 16408 2774 16436 4082
rect 16592 3058 16620 7142
rect 16776 6934 16804 7346
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 5409 16712 6734
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16776 6497 16804 6666
rect 16762 6488 16818 6497
rect 16762 6423 16818 6432
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16776 6089 16804 6190
rect 16762 6080 16818 6089
rect 16762 6015 16818 6024
rect 16670 5400 16726 5409
rect 16670 5335 16726 5344
rect 16684 5166 16712 5335
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 3670 16804 3878
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16868 3058 16896 9438
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16960 5302 16988 8502
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16316 2746 16436 2774
rect 12440 196 12492 202
rect 12440 138 12492 144
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16316 513 16344 2746
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 16684 1170 16712 2314
rect 16592 1142 16712 1170
rect 16592 800 16620 1142
rect 16960 800 16988 3606
rect 17052 2774 17080 9318
rect 17144 8974 17172 9318
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 7274 17172 8910
rect 17236 8430 17264 9472
rect 17592 9454 17644 9460
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17512 9042 17540 9318
rect 17408 9036 17460 9042
rect 17328 8996 17408 9024
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17236 6304 17264 8366
rect 17144 6276 17264 6304
rect 17144 5953 17172 6276
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17130 5944 17186 5953
rect 17130 5879 17186 5888
rect 17144 5370 17172 5879
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17144 3398 17172 4218
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17052 2746 17172 2774
rect 17144 2446 17172 2746
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17236 1494 17264 6054
rect 17328 4486 17356 8996
rect 17408 8978 17460 8984
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8566 17540 8842
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17420 8430 17448 8502
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17498 7984 17554 7993
rect 17498 7919 17554 7928
rect 17512 7886 17540 7919
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17420 7478 17448 7754
rect 17408 7472 17460 7478
rect 17460 7432 17540 7460
rect 17408 7414 17460 7420
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17420 5914 17448 7278
rect 17512 6934 17540 7432
rect 17604 7041 17632 7822
rect 17590 7032 17646 7041
rect 17590 6967 17646 6976
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17590 6896 17646 6905
rect 17590 6831 17646 6840
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17224 1488 17276 1494
rect 17224 1430 17276 1436
rect 17038 1320 17094 1329
rect 17038 1255 17094 1264
rect 17052 921 17080 1255
rect 17038 912 17094 921
rect 17038 847 17094 856
rect 17328 800 17356 3674
rect 17420 1193 17448 4966
rect 17512 1698 17540 6734
rect 17604 6662 17632 6831
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17604 5778 17632 6190
rect 17696 6186 17724 8298
rect 17788 6458 17816 9318
rect 17972 8906 18000 9676
rect 18340 9602 18368 9862
rect 18432 9654 18460 10610
rect 18524 10538 18552 10950
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18248 9574 18368 9602
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18248 9518 18276 9574
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18328 9512 18380 9518
rect 18380 9472 18460 9500
rect 18328 9454 18380 9460
rect 17960 8900 18012 8906
rect 17880 8860 17960 8888
rect 17880 8514 17908 8860
rect 17960 8842 18012 8848
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 17880 8486 18000 8514
rect 17972 7732 18000 8486
rect 17880 7704 18000 7732
rect 17880 7528 17908 7704
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17880 7500 18184 7528
rect 18156 7460 18184 7500
rect 18236 7472 18288 7478
rect 18156 7432 18236 7460
rect 18236 7414 18288 7420
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17684 6180 17736 6186
rect 17684 6122 17736 6128
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5302 17816 5510
rect 17776 5296 17828 5302
rect 17776 5238 17828 5244
rect 17880 5030 17908 7142
rect 18234 6896 18290 6905
rect 18234 6831 18290 6840
rect 18248 6730 18276 6831
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18340 6440 18368 8570
rect 18248 6412 18368 6440
rect 18248 6118 18276 6412
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18142 5944 18198 5953
rect 18142 5879 18198 5888
rect 18156 5710 18184 5879
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18328 5160 18380 5166
rect 18432 5137 18460 9472
rect 18510 8392 18566 8401
rect 18510 8327 18566 8336
rect 18524 6866 18552 8327
rect 18616 7342 18644 11154
rect 18694 11112 18750 11121
rect 18694 11047 18750 11056
rect 18708 10198 18736 11047
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18708 9926 18736 10134
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18694 9072 18750 9081
rect 18694 9007 18750 9016
rect 18708 8906 18736 9007
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18708 8401 18736 8434
rect 18694 8392 18750 8401
rect 18694 8327 18750 8336
rect 18800 8294 18828 15370
rect 18892 13530 18920 16238
rect 19076 15745 19104 17478
rect 19062 15736 19118 15745
rect 19062 15671 19118 15680
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19076 14074 19104 15506
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18892 7426 18920 12854
rect 18984 11354 19012 13874
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19076 12918 19104 13126
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18970 11248 19026 11257
rect 18970 11183 18972 11192
rect 19024 11183 19026 11192
rect 18972 11154 19024 11160
rect 18984 11082 19012 11154
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 19168 10713 19196 19722
rect 19260 18426 19288 20334
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19352 19514 19380 19722
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19352 18306 19380 19314
rect 19260 18278 19380 18306
rect 19260 15502 19288 18278
rect 19536 17678 19564 22374
rect 19628 21865 19656 22918
rect 19614 21856 19670 21865
rect 19614 21791 19670 21800
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19628 20942 19656 21626
rect 19720 21622 19748 23718
rect 19708 21616 19760 21622
rect 19708 21558 19760 21564
rect 19708 21072 19760 21078
rect 19708 21014 19760 21020
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19628 18766 19656 20198
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19720 16980 19748 21014
rect 19812 20058 19840 28070
rect 20076 28008 20128 28014
rect 20076 27950 20128 27956
rect 20088 27606 20116 27950
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 20180 27062 20208 28426
rect 20168 27056 20220 27062
rect 20168 26998 20220 27004
rect 20180 26790 20208 26998
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19904 23186 19932 24006
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19904 17252 19932 22918
rect 19996 18426 20024 24822
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 20088 22574 20116 23598
rect 20272 23118 20300 24346
rect 20364 24070 20392 29718
rect 20548 29306 20576 31622
rect 20640 30802 20668 32302
rect 20628 30796 20680 30802
rect 20628 30738 20680 30744
rect 20732 29646 20760 35430
rect 20824 33454 20852 35498
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 20812 33448 20864 33454
rect 20812 33390 20864 33396
rect 20916 33130 20944 33458
rect 20824 33102 20944 33130
rect 20824 32910 20852 33102
rect 20904 33040 20956 33046
rect 20904 32982 20956 32988
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20824 30598 20852 31962
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20916 29714 20944 32982
rect 21008 30326 21036 35430
rect 20996 30320 21048 30326
rect 20996 30262 21048 30268
rect 21100 29714 21128 38694
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21192 34678 21220 35566
rect 21180 34672 21232 34678
rect 21180 34614 21232 34620
rect 21192 34134 21220 34614
rect 21180 34128 21232 34134
rect 21180 34070 21232 34076
rect 21180 33924 21232 33930
rect 21180 33866 21232 33872
rect 21192 33522 21220 33866
rect 21180 33516 21232 33522
rect 21180 33458 21232 33464
rect 21180 30592 21232 30598
rect 21180 30534 21232 30540
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20444 28484 20496 28490
rect 20444 28426 20496 28432
rect 20456 27470 20484 28426
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20456 26450 20484 27406
rect 20444 26444 20496 26450
rect 20444 26386 20496 26392
rect 20640 26042 20668 29446
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20732 25498 20760 29106
rect 20824 28218 20852 29106
rect 21192 29102 21220 30534
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20904 28076 20956 28082
rect 20904 28018 20956 28024
rect 20916 27130 20944 28018
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 21100 27130 21128 27950
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26382 20852 26726
rect 21192 26518 21220 28562
rect 21284 28082 21312 41386
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 21364 34604 21416 34610
rect 21364 34546 21416 34552
rect 21376 33046 21404 34546
rect 21468 33862 21496 36110
rect 21744 35698 21772 46446
rect 21836 41414 21864 55186
rect 22388 53582 22416 55383
rect 22848 55214 22876 56222
rect 23032 56114 23060 56222
rect 23110 56200 23166 57000
rect 24122 56264 24178 56273
rect 23124 56114 23152 56200
rect 24122 56199 24178 56208
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 23032 56086 23152 56114
rect 22756 55186 22876 55214
rect 22376 53576 22428 53582
rect 22376 53518 22428 53524
rect 22100 53440 22152 53446
rect 22100 53382 22152 53388
rect 22112 49434 22140 53382
rect 22756 52494 22784 55186
rect 22834 54632 22890 54641
rect 22834 54567 22890 54576
rect 22848 53174 22876 54567
rect 23388 54052 23440 54058
rect 23388 53994 23440 54000
rect 23480 54052 23532 54058
rect 23480 53994 23532 54000
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23400 53825 23428 53994
rect 23386 53816 23442 53825
rect 23386 53751 23442 53760
rect 23296 53576 23348 53582
rect 23296 53518 23348 53524
rect 22836 53168 22888 53174
rect 22836 53110 22888 53116
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23308 52698 23336 53518
rect 23296 52692 23348 52698
rect 23296 52634 23348 52640
rect 23492 52494 23520 53994
rect 23940 53984 23992 53990
rect 23940 53926 23992 53932
rect 23756 53440 23808 53446
rect 23756 53382 23808 53388
rect 22744 52488 22796 52494
rect 22744 52430 22796 52436
rect 23480 52488 23532 52494
rect 23480 52430 23532 52436
rect 23768 52018 23796 53382
rect 23952 53106 23980 53926
rect 23940 53100 23992 53106
rect 23940 53042 23992 53048
rect 24136 52494 24164 56199
rect 24124 52488 24176 52494
rect 24124 52430 24176 52436
rect 23940 52352 23992 52358
rect 23940 52294 23992 52300
rect 23756 52012 23808 52018
rect 23756 51954 23808 51960
rect 22560 51808 22612 51814
rect 22560 51750 22612 51756
rect 22100 49428 22152 49434
rect 22100 49370 22152 49376
rect 22572 49230 22600 51750
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22560 49224 22612 49230
rect 22560 49166 22612 49172
rect 22652 49088 22704 49094
rect 22652 49030 22704 49036
rect 22664 47054 22692 49030
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22652 47048 22704 47054
rect 22652 46990 22704 46996
rect 22652 46368 22704 46374
rect 22652 46310 22704 46316
rect 22468 45824 22520 45830
rect 22468 45766 22520 45772
rect 22376 44736 22428 44742
rect 22376 44678 22428 44684
rect 21836 41386 21956 41414
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 21744 35222 21772 35634
rect 21732 35216 21784 35222
rect 21732 35158 21784 35164
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21456 33856 21508 33862
rect 21456 33798 21508 33804
rect 21652 33590 21680 34002
rect 21640 33584 21692 33590
rect 21640 33526 21692 33532
rect 21364 33040 21416 33046
rect 21364 32982 21416 32988
rect 21640 32768 21692 32774
rect 21640 32710 21692 32716
rect 21456 32496 21508 32502
rect 21456 32438 21508 32444
rect 21468 32026 21496 32438
rect 21652 32026 21680 32710
rect 21456 32020 21508 32026
rect 21456 31962 21508 31968
rect 21640 32020 21692 32026
rect 21640 31962 21692 31968
rect 21468 31482 21496 31962
rect 21744 31906 21772 35158
rect 21824 35012 21876 35018
rect 21824 34954 21876 34960
rect 21836 32609 21864 34954
rect 21822 32600 21878 32609
rect 21822 32535 21878 32544
rect 21652 31890 21864 31906
rect 21652 31884 21876 31890
rect 21652 31878 21824 31884
rect 21652 31822 21680 31878
rect 21824 31826 21876 31832
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21928 31754 21956 41386
rect 22192 37120 22244 37126
rect 22192 37062 22244 37068
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 22008 33856 22060 33862
rect 22008 33798 22060 33804
rect 22020 33658 22048 33798
rect 22008 33652 22060 33658
rect 22008 33594 22060 33600
rect 22112 33425 22140 34410
rect 22204 33930 22232 37062
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22296 36378 22324 36722
rect 22284 36372 22336 36378
rect 22284 36314 22336 36320
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22296 34082 22324 35226
rect 22388 35154 22416 44678
rect 22480 35834 22508 45766
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22664 35766 22692 46310
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 23480 43104 23532 43110
rect 23480 43046 23532 43052
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23492 40089 23520 43046
rect 23952 41478 23980 52294
rect 24136 51610 24164 52430
rect 24124 51604 24176 51610
rect 24124 51546 24176 51552
rect 24504 50386 24532 56200
rect 25320 54256 25372 54262
rect 25320 54198 25372 54204
rect 25228 54188 25280 54194
rect 25228 54130 25280 54136
rect 25136 54120 25188 54126
rect 25136 54062 25188 54068
rect 24584 53984 24636 53990
rect 24584 53926 24636 53932
rect 24596 53582 24624 53926
rect 24860 53712 24912 53718
rect 24860 53654 24912 53660
rect 24584 53576 24636 53582
rect 24584 53518 24636 53524
rect 24872 53174 24900 53654
rect 25148 53242 25176 54062
rect 25240 53786 25268 54130
rect 25228 53780 25280 53786
rect 25228 53722 25280 53728
rect 25136 53236 25188 53242
rect 25136 53178 25188 53184
rect 24860 53168 24912 53174
rect 24860 53110 24912 53116
rect 24582 53000 24638 53009
rect 24582 52935 24638 52944
rect 24596 52018 24624 52935
rect 24676 52896 24728 52902
rect 24676 52838 24728 52844
rect 24688 52494 24716 52838
rect 25332 52698 25360 54198
rect 25884 53718 25912 56200
rect 25872 53712 25924 53718
rect 25872 53654 25924 53660
rect 25320 52692 25372 52698
rect 25320 52634 25372 52640
rect 24676 52488 24728 52494
rect 24676 52430 24728 52436
rect 24950 52184 25006 52193
rect 24950 52119 25006 52128
rect 24964 52086 24992 52119
rect 24952 52080 25004 52086
rect 24952 52022 25004 52028
rect 24584 52012 24636 52018
rect 24584 51954 24636 51960
rect 24596 51610 24624 51954
rect 24584 51604 24636 51610
rect 24584 51546 24636 51552
rect 24964 51542 24992 52022
rect 24952 51536 25004 51542
rect 24952 51478 25004 51484
rect 24950 51368 25006 51377
rect 24950 51303 24952 51312
rect 25004 51303 25006 51312
rect 24952 51274 25004 51280
rect 25044 51264 25096 51270
rect 25044 51206 25096 51212
rect 24952 50924 25004 50930
rect 24952 50866 25004 50872
rect 24584 50720 24636 50726
rect 24584 50662 24636 50668
rect 24596 50522 24624 50662
rect 24964 50561 24992 50866
rect 24950 50552 25006 50561
rect 24584 50516 24636 50522
rect 24950 50487 25006 50496
rect 24584 50458 24636 50464
rect 24492 50380 24544 50386
rect 24492 50322 24544 50328
rect 24768 49768 24820 49774
rect 24768 49710 24820 49716
rect 24780 47705 24808 49710
rect 24860 48000 24912 48006
rect 24860 47942 24912 47948
rect 24766 47696 24822 47705
rect 24766 47631 24822 47640
rect 24872 47025 24900 47942
rect 24858 47016 24914 47025
rect 24858 46951 24914 46960
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 44033 24808 44338
rect 25056 44198 25084 51206
rect 25504 50176 25556 50182
rect 25504 50118 25556 50124
rect 25516 49842 25544 50118
rect 25504 49836 25556 49842
rect 25504 49778 25556 49784
rect 25516 49745 25544 49778
rect 25502 49736 25558 49745
rect 25502 49671 25558 49680
rect 25136 49156 25188 49162
rect 25136 49098 25188 49104
rect 25148 48929 25176 49098
rect 25228 49088 25280 49094
rect 25228 49030 25280 49036
rect 25134 48920 25190 48929
rect 25134 48855 25190 48864
rect 25136 48544 25188 48550
rect 25136 48486 25188 48492
rect 25148 48142 25176 48486
rect 25136 48136 25188 48142
rect 25134 48104 25136 48113
rect 25188 48104 25190 48113
rect 25134 48039 25190 48048
rect 25240 47569 25268 49030
rect 25320 47660 25372 47666
rect 25320 47602 25372 47608
rect 25226 47560 25282 47569
rect 25226 47495 25282 47504
rect 25332 47297 25360 47602
rect 25780 47456 25832 47462
rect 25780 47398 25832 47404
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25332 46578 25360 46854
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25320 45280 25372 45286
rect 25320 45222 25372 45228
rect 25332 44878 25360 45222
rect 25320 44872 25372 44878
rect 25318 44840 25320 44849
rect 25372 44840 25374 44849
rect 25318 44775 25374 44784
rect 25044 44192 25096 44198
rect 25044 44134 25096 44140
rect 24766 44024 24822 44033
rect 24766 43959 24822 43968
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25516 43382 25544 43590
rect 25504 43376 25556 43382
rect 25504 43318 25556 43324
rect 25516 43217 25544 43318
rect 25502 43208 25558 43217
rect 25502 43143 25558 43152
rect 25226 42664 25282 42673
rect 25136 42628 25188 42634
rect 25226 42599 25282 42608
rect 25136 42570 25188 42576
rect 25148 42401 25176 42570
rect 25240 42566 25268 42599
rect 25228 42560 25280 42566
rect 25228 42502 25280 42508
rect 25134 42392 25190 42401
rect 25134 42327 25190 42336
rect 25320 42016 25372 42022
rect 25320 41958 25372 41964
rect 24858 41576 24914 41585
rect 24858 41511 24914 41520
rect 25134 41576 25190 41585
rect 25134 41511 25136 41520
rect 24872 41478 24900 41511
rect 25188 41511 25190 41520
rect 25136 41482 25188 41488
rect 23940 41472 23992 41478
rect 23940 41414 23992 41420
rect 24860 41472 24912 41478
rect 24860 41414 24912 41420
rect 25332 41138 25360 41958
rect 24860 41132 24912 41138
rect 24860 41074 24912 41080
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 23848 40928 23900 40934
rect 23848 40870 23900 40876
rect 23478 40080 23534 40089
rect 23478 40015 23534 40024
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22744 38208 22796 38214
rect 22744 38150 22796 38156
rect 22652 35760 22704 35766
rect 22652 35702 22704 35708
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 22376 35148 22428 35154
rect 22376 35090 22428 35096
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22480 34354 22508 34886
rect 22572 34474 22600 35566
rect 22652 35216 22704 35222
rect 22652 35158 22704 35164
rect 22664 34626 22692 35158
rect 22756 35057 22784 38150
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23480 37664 23532 37670
rect 23480 37606 23532 37612
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23492 37262 23520 37606
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23204 36032 23256 36038
rect 23204 35974 23256 35980
rect 23216 35698 23244 35974
rect 23204 35692 23256 35698
rect 23204 35634 23256 35640
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23308 35154 23336 36110
rect 23400 35698 23428 36518
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 22742 35048 22798 35057
rect 22742 34983 22798 34992
rect 22664 34598 22784 34626
rect 22652 34536 22704 34542
rect 22652 34478 22704 34484
rect 22560 34468 22612 34474
rect 22560 34410 22612 34416
rect 22480 34326 22600 34354
rect 22296 34054 22416 34082
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22098 33416 22154 33425
rect 22098 33351 22154 33360
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 22020 32910 22048 33254
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 21744 31726 21956 31754
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21284 27130 21312 28018
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20718 25392 20774 25401
rect 20718 25327 20774 25336
rect 20996 25356 21048 25362
rect 20732 25294 20760 25327
rect 20996 25298 21048 25304
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20732 24954 20760 25230
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20904 25152 20956 25158
rect 20904 25094 20956 25100
rect 20824 24993 20852 25094
rect 20810 24984 20866 24993
rect 20720 24948 20772 24954
rect 20810 24919 20866 24928
rect 20720 24890 20772 24896
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 20352 24064 20404 24070
rect 20456 24041 20484 24074
rect 20352 24006 20404 24012
rect 20442 24032 20498 24041
rect 20442 23967 20498 23976
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20640 23118 20668 23462
rect 20732 23186 20760 24142
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 20180 22506 20208 23054
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 22642 20760 22918
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20180 21554 20208 22170
rect 20824 22030 20852 23122
rect 20916 22778 20944 25094
rect 21008 24274 21036 25298
rect 21192 25226 21220 26454
rect 21284 26042 21312 26862
rect 21376 26450 21404 31146
rect 21468 29646 21496 31418
rect 21744 30274 21772 31726
rect 22020 31634 22048 32846
rect 22112 31793 22140 33050
rect 22296 32978 22324 33526
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22296 32502 22324 32914
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22098 31784 22154 31793
rect 22098 31719 22154 31728
rect 22020 31606 22140 31634
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22020 30938 22048 31282
rect 22112 31249 22140 31606
rect 22098 31240 22154 31249
rect 22098 31175 22154 31184
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 21824 30660 21876 30666
rect 21824 30602 21876 30608
rect 21836 30394 21864 30602
rect 21824 30388 21876 30394
rect 21824 30330 21876 30336
rect 22284 30388 22336 30394
rect 22284 30330 22336 30336
rect 21560 30246 21772 30274
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21364 26444 21416 26450
rect 21364 26386 21416 26392
rect 21560 26042 21588 30246
rect 21732 30116 21784 30122
rect 21732 30058 21784 30064
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21548 26036 21600 26042
rect 21548 25978 21600 25984
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21180 25220 21232 25226
rect 21180 25162 21232 25168
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21284 24614 21312 24754
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 21008 23610 21036 24210
rect 21284 24138 21312 24550
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21008 23582 21220 23610
rect 21088 23520 21140 23526
rect 20994 23488 21050 23497
rect 21088 23462 21140 23468
rect 20994 23423 21050 23432
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20824 21690 20852 21830
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20088 19446 20116 19858
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20088 19174 20116 19382
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20272 18970 20300 21490
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20364 19718 20392 20946
rect 20456 20806 20484 21490
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20824 20806 20852 21422
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20628 20800 20680 20806
rect 20812 20800 20864 20806
rect 20628 20742 20680 20748
rect 20810 20768 20812 20777
rect 20864 20768 20866 20777
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20180 18086 20208 18566
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20364 17762 20392 19654
rect 20272 17734 20392 17762
rect 19904 17224 20024 17252
rect 19444 16952 19748 16980
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19352 14074 19380 15982
rect 19444 14074 19472 16952
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19720 16590 19748 16730
rect 19708 16584 19760 16590
rect 19628 16544 19708 16572
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19536 15337 19564 15370
rect 19522 15328 19578 15337
rect 19522 15263 19578 15272
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19352 13682 19380 14010
rect 19536 14006 19564 14350
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19352 13654 19564 13682
rect 19338 13560 19394 13569
rect 19338 13495 19340 13504
rect 19392 13495 19394 13504
rect 19340 13466 19392 13472
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19260 12986 19288 13262
rect 19352 13190 19380 13466
rect 19536 13394 19564 13654
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19444 12986 19472 13330
rect 19536 13161 19564 13330
rect 19522 13152 19578 13161
rect 19522 13087 19578 13096
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19628 12918 19656 16544
rect 19708 16526 19760 16532
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19352 12434 19380 12854
rect 19352 12406 19472 12434
rect 19444 12102 19472 12406
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11830 19472 12038
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19338 11384 19394 11393
rect 19338 11319 19340 11328
rect 19392 11319 19394 11328
rect 19340 11290 19392 11296
rect 19154 10704 19210 10713
rect 19210 10662 19288 10690
rect 19154 10639 19210 10648
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 9586 19012 9862
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18984 8430 19012 9318
rect 19168 9110 19196 10542
rect 19260 10130 19288 10662
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18800 7398 18920 7426
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18604 6860 18656 6866
rect 18656 6820 18736 6848
rect 18604 6802 18656 6808
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18328 5102 18380 5108
rect 18418 5128 18474 5137
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17604 3398 17632 4014
rect 17788 3641 17816 4762
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17774 3632 17830 3641
rect 17774 3567 17830 3576
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17500 1692 17552 1698
rect 17500 1634 17552 1640
rect 17406 1184 17462 1193
rect 17406 1119 17462 1128
rect 17696 800 17724 2586
rect 17880 2417 17908 4626
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 18064 3602 18092 3975
rect 18340 3738 18368 5102
rect 18418 5063 18474 5072
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18432 3670 18460 4490
rect 18524 4214 18552 6598
rect 18708 5846 18736 6820
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18512 4208 18564 4214
rect 18512 4150 18564 4156
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18524 2961 18552 4014
rect 18510 2952 18566 2961
rect 18510 2887 18566 2896
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17866 2408 17922 2417
rect 18248 2394 18276 2790
rect 18616 2666 18644 4966
rect 18800 4282 18828 7398
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18432 2638 18644 2666
rect 18248 2366 18368 2394
rect 17866 2343 17922 2352
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 16302 504 16358 513
rect 16302 439 16358 448
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2366
rect 18432 800 18460 2638
rect 18708 921 18736 3470
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18694 912 18750 921
rect 18694 847 18750 856
rect 18800 800 18828 3130
rect 18892 3058 18920 7278
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18878 2952 18934 2961
rect 18878 2887 18934 2896
rect 18892 1154 18920 2887
rect 18984 2514 19012 8230
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19076 2650 19104 7754
rect 19168 2961 19196 9046
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8566 19288 8774
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19260 8430 19288 8502
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19352 8294 19380 10610
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19352 7750 19380 7958
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19260 7562 19288 7686
rect 19260 7534 19380 7562
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 6390 19288 7346
rect 19352 7177 19380 7534
rect 19338 7168 19394 7177
rect 19338 7103 19394 7112
rect 19248 6384 19300 6390
rect 19300 6344 19380 6372
rect 19248 6326 19300 6332
rect 19352 5953 19380 6344
rect 19338 5944 19394 5953
rect 19248 5908 19300 5914
rect 19338 5879 19394 5888
rect 19248 5850 19300 5856
rect 19260 5001 19288 5850
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19246 4992 19302 5001
rect 19246 4927 19302 4936
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19260 4282 19288 4490
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19154 2952 19210 2961
rect 19154 2887 19210 2896
rect 19352 2774 19380 5714
rect 19444 4622 19472 9862
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19430 4176 19486 4185
rect 19430 4111 19486 4120
rect 19168 2746 19380 2774
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 18880 1148 18932 1154
rect 18880 1090 18932 1096
rect 19168 800 19196 2746
rect 19444 2446 19472 4111
rect 19536 4026 19564 12174
rect 19720 11529 19748 15370
rect 19798 14784 19854 14793
rect 19798 14719 19854 14728
rect 19812 12918 19840 14719
rect 19800 12912 19852 12918
rect 19800 12854 19852 12860
rect 19812 12442 19840 12854
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19706 11520 19762 11529
rect 19706 11455 19762 11464
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19720 10266 19748 10474
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19628 8838 19656 9454
rect 19812 9330 19840 11222
rect 19904 9654 19932 15370
rect 19996 12434 20024 17224
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20088 15094 20116 15302
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20088 14482 20116 15030
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19996 12406 20116 12434
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19996 10266 20024 12106
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19996 9489 20024 9590
rect 19982 9480 20038 9489
rect 19982 9415 20038 9424
rect 19720 9302 19840 9330
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19628 7993 19656 8026
rect 19614 7984 19670 7993
rect 19614 7919 19670 7928
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19628 7410 19656 7754
rect 19720 7750 19748 9302
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19812 7818 19840 9114
rect 20088 7970 20116 12406
rect 20272 12374 20300 17734
rect 20456 15910 20484 20334
rect 20640 20262 20668 20742
rect 20810 20703 20866 20712
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20640 19689 20668 19926
rect 20732 19825 20760 20402
rect 20810 19952 20866 19961
rect 20810 19887 20866 19896
rect 20824 19854 20852 19887
rect 20812 19848 20864 19854
rect 20718 19816 20774 19825
rect 20812 19790 20864 19796
rect 20718 19751 20774 19760
rect 20626 19680 20682 19689
rect 20626 19615 20682 19624
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18902 20576 19110
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20350 15056 20406 15065
rect 20350 14991 20406 15000
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20180 11830 20208 12174
rect 20272 12102 20300 12310
rect 20364 12238 20392 14991
rect 20442 13968 20498 13977
rect 20442 13903 20444 13912
rect 20496 13903 20498 13912
rect 20444 13874 20496 13880
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12306 20484 12718
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20548 11914 20576 18838
rect 20640 16658 20668 19450
rect 20810 18728 20866 18737
rect 20810 18663 20866 18672
rect 20824 16794 20852 18663
rect 20916 18630 20944 21286
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 21008 17882 21036 23423
rect 21100 22234 21128 23462
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 21100 22030 21128 22170
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21192 21894 21220 23582
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21100 21622 21128 21830
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 21192 20754 21220 21830
rect 21284 20913 21312 23462
rect 21376 22778 21404 24686
rect 21468 23730 21496 25230
rect 21560 24410 21588 25842
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 21652 24206 21680 26726
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21456 23588 21508 23594
rect 21456 23530 21508 23536
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21468 22098 21496 23530
rect 21548 23316 21600 23322
rect 21548 23258 21600 23264
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21270 20904 21326 20913
rect 21270 20839 21326 20848
rect 21192 20726 21312 20754
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 21100 16980 21128 20198
rect 21284 17202 21312 20726
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21100 16952 21220 16980
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20640 15570 20668 16594
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15162 20668 15506
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20640 14958 20668 15098
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20732 14890 20760 16390
rect 20824 16182 20852 16730
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 13870 20668 14758
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20626 13424 20682 13433
rect 20626 13359 20628 13368
rect 20680 13359 20682 13368
rect 20628 13330 20680 13336
rect 20718 13288 20774 13297
rect 20718 13223 20774 13232
rect 20732 13190 20760 13223
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20272 11886 20576 11914
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20272 11762 20300 11886
rect 20352 11824 20404 11830
rect 20640 11778 20668 12922
rect 20720 12640 20772 12646
rect 20718 12608 20720 12617
rect 20772 12608 20774 12617
rect 20718 12543 20774 12552
rect 20352 11766 20404 11772
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20364 11558 20392 11766
rect 20456 11750 20668 11778
rect 20824 11762 20852 15846
rect 20996 15360 21048 15366
rect 20902 15328 20958 15337
rect 20996 15302 21048 15308
rect 20902 15263 20958 15272
rect 20916 15094 20944 15263
rect 21008 15162 21036 15302
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 20916 14414 20944 14826
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13870 20944 14214
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20916 12442 20944 13806
rect 21100 13530 21128 16050
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21192 13326 21220 16952
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 16046 21312 16390
rect 21376 16250 21404 21626
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21468 20806 21496 21558
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21560 20602 21588 23258
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21560 20466 21588 20538
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17202 21496 17614
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21560 16590 21588 20198
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21652 16454 21680 23190
rect 21744 22710 21772 30058
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21928 28490 21956 29582
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 22006 29064 22062 29073
rect 22006 28999 22008 29008
rect 22060 28999 22062 29008
rect 22008 28970 22060 28976
rect 22112 28642 22140 29514
rect 22020 28614 22140 28642
rect 21916 28484 21968 28490
rect 21916 28426 21968 28432
rect 22020 28082 22048 28614
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21928 27606 21956 27814
rect 21916 27600 21968 27606
rect 21916 27542 21968 27548
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21836 24993 21864 27066
rect 22020 26994 22048 28018
rect 22100 27124 22152 27130
rect 22100 27066 22152 27072
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22020 26450 22048 26930
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 21928 26330 21956 26386
rect 21928 26314 22048 26330
rect 21928 26308 22060 26314
rect 21928 26302 22008 26308
rect 22008 26250 22060 26256
rect 22112 26246 22140 27066
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 21916 25492 21968 25498
rect 21916 25434 21968 25440
rect 21928 25294 21956 25434
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21916 25152 21968 25158
rect 22112 25140 22140 25978
rect 21968 25112 22140 25140
rect 21916 25094 21968 25100
rect 21822 24984 21878 24993
rect 21822 24919 21878 24928
rect 21916 24880 21968 24886
rect 21836 24840 21916 24868
rect 21836 23730 21864 24840
rect 21916 24822 21968 24828
rect 22112 24614 22140 25112
rect 22204 24682 22232 28358
rect 22296 28150 22324 30330
rect 22388 28762 22416 34054
rect 22572 32314 22600 34326
rect 22480 32286 22600 32314
rect 22480 29306 22508 32286
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22572 31890 22600 32166
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22664 30734 22692 34478
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22756 30274 22784 34598
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22848 32994 22876 34546
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23308 33114 23336 35090
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23400 34950 23428 35022
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23400 34490 23428 34886
rect 23400 34462 23520 34490
rect 23388 34400 23440 34406
rect 23388 34342 23440 34348
rect 23400 34134 23428 34342
rect 23388 34128 23440 34134
rect 23388 34070 23440 34076
rect 23492 33946 23520 34462
rect 23400 33918 23520 33946
rect 23204 33108 23256 33114
rect 23204 33050 23256 33056
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 22848 32978 22968 32994
rect 22848 32972 22980 32978
rect 22848 32966 22928 32972
rect 22848 30938 22876 32966
rect 22928 32914 22980 32920
rect 23020 32836 23072 32842
rect 23020 32778 23072 32784
rect 23032 32502 23060 32778
rect 23216 32774 23244 33050
rect 23400 32994 23428 33918
rect 23676 33318 23704 37810
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23308 32966 23428 32994
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 23216 31482 23244 31758
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22836 30796 22888 30802
rect 22836 30738 22888 30744
rect 22664 30246 22784 30274
rect 22560 30116 22612 30122
rect 22560 30058 22612 30064
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22480 28558 22508 28902
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 22284 28144 22336 28150
rect 22284 28086 22336 28092
rect 22296 27588 22324 28086
rect 22296 27560 22508 27588
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 26897 22324 27270
rect 22480 27130 22508 27560
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22376 27056 22428 27062
rect 22376 26998 22428 27004
rect 22282 26888 22338 26897
rect 22282 26823 22338 26832
rect 22388 26081 22416 26998
rect 22466 26752 22522 26761
rect 22466 26687 22522 26696
rect 22374 26072 22430 26081
rect 22374 26007 22430 26016
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21836 23322 21864 23666
rect 21928 23594 21956 24142
rect 22006 23624 22062 23633
rect 21916 23588 21968 23594
rect 22006 23559 22062 23568
rect 21916 23530 21968 23536
rect 22020 23526 22048 23559
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 22112 23338 22140 24550
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 22020 23310 22140 23338
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21732 22704 21784 22710
rect 21732 22646 21784 22652
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21744 19786 21772 22034
rect 21836 21078 21864 23054
rect 22020 22522 22048 23310
rect 22098 23216 22154 23225
rect 22098 23151 22154 23160
rect 22112 22642 22140 23151
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22020 22494 22232 22522
rect 21914 22128 21970 22137
rect 21914 22063 21970 22072
rect 21928 21865 21956 22063
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 21914 21856 21970 21865
rect 21914 21791 21970 21800
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21824 20936 21876 20942
rect 21822 20904 21824 20913
rect 21876 20904 21878 20913
rect 21822 20839 21878 20848
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21732 19780 21784 19786
rect 21732 19722 21784 19728
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 14929 21680 15982
rect 21836 15978 21864 20742
rect 21928 18970 21956 21791
rect 22020 21729 22048 21898
rect 22006 21720 22062 21729
rect 22006 21655 22062 21664
rect 22204 21622 22232 22494
rect 22192 21616 22244 21622
rect 22190 21584 22192 21593
rect 22244 21584 22246 21593
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22100 21548 22152 21554
rect 22296 21554 22324 24074
rect 22190 21519 22246 21528
rect 22284 21548 22336 21554
rect 22100 21490 22152 21496
rect 22284 21490 22336 21496
rect 22020 21078 22048 21490
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 22006 20360 22062 20369
rect 22006 20295 22008 20304
rect 22060 20295 22062 20304
rect 22008 20266 22060 20272
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 22112 18426 22140 21490
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22296 20398 22324 21354
rect 22388 20602 22416 24550
rect 22480 21622 22508 26687
rect 22572 25294 22600 30058
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22468 21480 22520 21486
rect 22466 21448 22468 21457
rect 22520 21448 22522 21457
rect 22466 21383 22522 21392
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22204 18698 22232 19790
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22296 18834 22324 19450
rect 22388 19446 22416 19654
rect 22376 19440 22428 19446
rect 22376 19382 22428 19388
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22284 18692 22336 18698
rect 22284 18634 22336 18640
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 21914 18320 21970 18329
rect 21914 18255 21970 18264
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21836 15570 21864 15914
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21638 14920 21694 14929
rect 21638 14855 21694 14864
rect 21652 14822 21680 14855
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21270 14376 21326 14385
rect 21270 14311 21326 14320
rect 21284 13734 21312 14311
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20994 12472 21050 12481
rect 20904 12436 20956 12442
rect 20994 12407 21050 12416
rect 20904 12378 20956 12384
rect 21008 11762 21036 12407
rect 20812 11756 20864 11762
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20166 11248 20222 11257
rect 20272 11218 20300 11494
rect 20166 11183 20168 11192
rect 20220 11183 20222 11192
rect 20260 11212 20312 11218
rect 20168 11154 20220 11160
rect 20260 11154 20312 11160
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20180 9874 20208 10950
rect 20272 10742 20300 10950
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20364 10674 20392 11018
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20258 9888 20314 9897
rect 20180 9846 20258 9874
rect 20258 9823 20314 9832
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19904 7954 20116 7970
rect 19892 7948 20116 7954
rect 19944 7942 20116 7948
rect 19892 7890 19944 7896
rect 19800 7812 19852 7818
rect 19800 7754 19852 7760
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19616 7200 19668 7206
rect 19904 7177 19932 7686
rect 19616 7142 19668 7148
rect 19890 7168 19946 7177
rect 19628 7002 19656 7142
rect 19890 7103 19946 7112
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19628 6440 19656 6938
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19892 6928 19944 6934
rect 19892 6870 19944 6876
rect 19812 6798 19840 6870
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19628 6412 19748 6440
rect 19720 6186 19748 6412
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19616 6112 19668 6118
rect 19614 6080 19616 6089
rect 19668 6080 19670 6089
rect 19614 6015 19670 6024
rect 19706 5944 19762 5953
rect 19706 5879 19762 5888
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19628 5370 19656 5646
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19720 4758 19748 5879
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 19720 4162 19748 4694
rect 19628 4146 19748 4162
rect 19616 4140 19748 4146
rect 19668 4134 19748 4140
rect 19616 4082 19668 4088
rect 19708 4072 19760 4078
rect 19706 4040 19708 4049
rect 19760 4040 19762 4049
rect 19536 3998 19656 4026
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19536 800 19564 2926
rect 19628 1018 19656 3998
rect 19706 3975 19762 3984
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19720 3602 19748 3878
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19616 1012 19668 1018
rect 19616 954 19668 960
rect 19720 882 19748 3402
rect 19812 1970 19840 5102
rect 19904 4826 19932 6870
rect 19996 5642 20024 7754
rect 20088 6866 20116 7942
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20074 6760 20130 6769
rect 20074 6695 20076 6704
rect 20128 6695 20130 6704
rect 20076 6666 20128 6672
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19982 5128 20038 5137
rect 19982 5063 20038 5072
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 19904 3913 19932 4150
rect 19996 3942 20024 5063
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 3936 20036 3942
rect 19890 3904 19946 3913
rect 19984 3878 20036 3884
rect 19890 3839 19946 3848
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19800 1964 19852 1970
rect 19800 1906 19852 1912
rect 19708 876 19760 882
rect 19708 818 19760 824
rect 19904 800 19932 2790
rect 20088 1222 20116 4558
rect 20180 3942 20208 8434
rect 20272 8362 20300 9823
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20258 7984 20314 7993
rect 20258 7919 20260 7928
rect 20312 7919 20314 7928
rect 20260 7890 20312 7896
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20272 6118 20300 6258
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20272 5914 20300 6054
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 20272 800 20300 4082
rect 20364 4078 20392 9522
rect 20456 8634 20484 11750
rect 20812 11698 20864 11704
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20640 10062 20668 11630
rect 21100 11354 21128 13126
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 8090 20484 8230
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20456 5574 20484 6394
rect 20548 6118 20576 9658
rect 20640 9042 20668 9998
rect 20732 9722 20760 10202
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20626 8528 20682 8537
rect 20626 8463 20682 8472
rect 20640 6118 20668 8463
rect 20718 7848 20774 7857
rect 20718 7783 20774 7792
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20732 6066 20760 7783
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20824 6225 20852 6734
rect 20810 6216 20866 6225
rect 20810 6151 20866 6160
rect 20732 6038 20852 6066
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20456 4690 20484 5510
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20364 2009 20392 3878
rect 20456 3602 20484 4626
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20548 2774 20576 5714
rect 20824 5710 20852 6038
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20732 4729 20760 5578
rect 20718 4720 20774 4729
rect 20718 4655 20774 4664
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4554 20852 4626
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20916 4162 20944 10202
rect 21100 9625 21128 10610
rect 21086 9616 21142 9625
rect 21086 9551 21142 9560
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 20732 4134 20944 4162
rect 20732 4078 20760 4134
rect 20720 4072 20772 4078
rect 20626 4040 20682 4049
rect 20720 4014 20772 4020
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20626 3975 20682 3984
rect 20640 3058 20668 3975
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20732 3194 20760 3538
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20548 2746 20668 2774
rect 20350 2000 20406 2009
rect 20350 1935 20406 1944
rect 20640 800 20668 2746
rect 20824 1057 20852 4014
rect 21008 2530 21036 9386
rect 21284 8514 21312 12582
rect 21376 11898 21404 13194
rect 21454 12744 21510 12753
rect 21454 12679 21510 12688
rect 21468 12646 21496 12679
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21560 9450 21588 14758
rect 21730 14648 21786 14657
rect 21730 14583 21786 14592
rect 21744 14550 21772 14583
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21652 12646 21680 14418
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21744 11830 21772 13738
rect 21836 12866 21864 13874
rect 21928 13326 21956 18255
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 22020 17202 22048 18090
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22020 14482 22048 14894
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22006 14376 22062 14385
rect 22006 14311 22008 14320
rect 22060 14311 22062 14320
rect 22008 14282 22060 14288
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21928 12986 21956 13262
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22020 12918 22048 14282
rect 22112 14006 22140 18022
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22204 16794 22232 17206
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22098 13016 22154 13025
rect 22098 12951 22154 12960
rect 22008 12912 22060 12918
rect 21836 12838 21956 12866
rect 22008 12854 22060 12860
rect 22112 12850 22140 12951
rect 21928 12782 21956 12838
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21638 11112 21694 11121
rect 21638 11047 21640 11056
rect 21692 11047 21694 11056
rect 21640 11018 21692 11024
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21548 8560 21600 8566
rect 21284 8486 21404 8514
rect 21548 8502 21600 8508
rect 21180 8424 21232 8430
rect 21232 8384 21312 8412
rect 21180 8366 21232 8372
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21192 4865 21220 5170
rect 21178 4856 21234 4865
rect 21178 4791 21234 4800
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 20916 2502 21036 2530
rect 20810 1048 20866 1057
rect 20810 983 20866 992
rect 20916 950 20944 2502
rect 21100 2394 21128 4626
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 21192 3534 21220 4490
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21284 3058 21312 8384
rect 21376 4214 21404 8486
rect 21560 5250 21588 8502
rect 21652 5914 21680 11018
rect 21730 9616 21786 9625
rect 21730 9551 21786 9560
rect 21744 6458 21772 9551
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21560 5222 21680 5250
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 21560 4146 21588 5102
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 21008 2366 21128 2394
rect 20904 944 20956 950
rect 20904 886 20956 892
rect 21008 800 21036 2366
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21100 1086 21128 2246
rect 21284 1290 21312 2246
rect 21272 1284 21324 1290
rect 21272 1226 21324 1232
rect 21088 1080 21140 1086
rect 21088 1022 21140 1028
rect 21376 800 21404 3946
rect 21468 2990 21496 4014
rect 21652 3942 21680 5222
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21652 1873 21680 3470
rect 21638 1864 21694 1873
rect 21638 1799 21694 1808
rect 21744 800 21772 6190
rect 21836 2446 21864 12718
rect 21928 10810 21956 12718
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 22020 10062 22048 12106
rect 22008 10056 22060 10062
rect 21928 10016 22008 10044
rect 21928 8974 21956 10016
rect 22008 9998 22060 10004
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22098 8936 22154 8945
rect 22020 7410 22048 8910
rect 22098 8871 22100 8880
rect 22152 8871 22154 8880
rect 22100 8842 22152 8848
rect 22098 7440 22154 7449
rect 22008 7404 22060 7410
rect 22098 7375 22154 7384
rect 22008 7346 22060 7352
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21928 3346 21956 6666
rect 22020 5574 22048 7346
rect 22112 7206 22140 7375
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22098 6352 22154 6361
rect 22098 6287 22100 6296
rect 22152 6287 22154 6296
rect 22100 6258 22152 6264
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22112 4570 22140 5306
rect 22020 4542 22140 4570
rect 22020 3466 22048 4542
rect 22204 4146 22232 14214
rect 22296 11014 22324 18634
rect 22388 18630 22416 19382
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22388 18358 22416 18566
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22388 15094 22416 18294
rect 22572 17678 22600 25094
rect 22664 24750 22692 30246
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22756 29578 22784 30126
rect 22848 29782 22876 30738
rect 23308 30161 23336 32966
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23400 31346 23428 32370
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23294 30152 23350 30161
rect 23294 30087 23350 30096
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22744 29572 22796 29578
rect 22744 29514 22796 29520
rect 23400 29345 23428 29786
rect 23386 29336 23442 29345
rect 23386 29271 23442 29280
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 22744 28008 22796 28014
rect 22744 27950 22796 27956
rect 22756 25106 22784 27950
rect 22848 27588 22876 29106
rect 23388 29096 23440 29102
rect 23202 29064 23258 29073
rect 23492 29050 23520 33254
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23584 29170 23612 29446
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23440 29044 23520 29050
rect 23388 29038 23520 29044
rect 23202 28999 23204 29008
rect 23256 28999 23258 29008
rect 23296 29028 23348 29034
rect 23204 28970 23256 28976
rect 23400 29022 23520 29038
rect 23296 28970 23348 28976
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23020 28688 23072 28694
rect 23020 28630 23072 28636
rect 23032 27878 23060 28630
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23308 27674 23336 28970
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23584 27878 23612 28494
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23400 27713 23428 27814
rect 23386 27704 23442 27713
rect 23296 27668 23348 27674
rect 23386 27639 23442 27648
rect 23480 27668 23532 27674
rect 23296 27610 23348 27616
rect 23480 27610 23532 27616
rect 22848 27560 22968 27588
rect 22834 27432 22890 27441
rect 22940 27402 22968 27560
rect 23492 27554 23520 27610
rect 23400 27526 23520 27554
rect 22834 27367 22890 27376
rect 22928 27396 22980 27402
rect 22848 27334 22876 27367
rect 22928 27338 22980 27344
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22940 27146 22968 27338
rect 22848 27118 22968 27146
rect 22848 25226 22876 27118
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23296 26444 23348 26450
rect 23296 26386 23348 26392
rect 23308 25974 23336 26386
rect 23400 26058 23428 27526
rect 23400 26030 23520 26058
rect 23296 25968 23348 25974
rect 23388 25968 23440 25974
rect 23296 25910 23348 25916
rect 23386 25936 23388 25945
rect 23440 25936 23442 25945
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22756 25078 22876 25106
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 20534 22692 23598
rect 22742 21720 22798 21729
rect 22742 21655 22798 21664
rect 22652 20528 22704 20534
rect 22652 20470 22704 20476
rect 22756 19938 22784 21655
rect 22848 20058 22876 25078
rect 23308 24750 23336 25910
rect 23386 25871 23442 25880
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24290 23336 24686
rect 23216 24262 23336 24290
rect 23216 23662 23244 24262
rect 23400 23798 23428 25774
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23204 23656 23256 23662
rect 23492 23610 23520 26030
rect 23204 23598 23256 23604
rect 23400 23582 23520 23610
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23400 23050 23428 23582
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 21480 23256 21486
rect 23256 21428 23336 21434
rect 23204 21422 23336 21428
rect 23216 21406 23336 21422
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23124 20262 23152 20810
rect 23202 20768 23258 20777
rect 23202 20703 23258 20712
rect 23216 20602 23244 20703
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 23308 20466 23336 21406
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22756 19910 22876 19938
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22466 17096 22522 17105
rect 22466 17031 22468 17040
rect 22520 17031 22522 17040
rect 22468 17002 22520 17008
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22572 13190 22600 14554
rect 22664 13530 22692 17614
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22388 10742 22416 12854
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22376 10736 22428 10742
rect 22296 10696 22376 10724
rect 22296 10606 22324 10696
rect 22376 10678 22428 10684
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22296 9926 22324 10542
rect 22376 10532 22428 10538
rect 22376 10474 22428 10480
rect 22388 10198 22416 10474
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 21928 3318 22232 3346
rect 22098 3088 22154 3097
rect 22098 3023 22100 3032
rect 22152 3023 22154 3032
rect 22100 2994 22152 3000
rect 22204 2774 22232 3318
rect 22296 3233 22324 9454
rect 22480 9382 22508 12310
rect 22664 12306 22692 12718
rect 22756 12442 22784 19246
rect 22848 18086 22876 19910
rect 23308 19514 23336 20402
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23400 19553 23428 19722
rect 23386 19544 23442 19553
rect 23296 19508 23348 19514
rect 23386 19479 23442 19488
rect 23296 19450 23348 19456
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23308 18290 23336 19450
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23386 18184 23442 18193
rect 23492 18154 23520 19178
rect 23584 18834 23612 27814
rect 23676 27130 23704 30126
rect 23768 29646 23796 34478
rect 23860 33658 23888 40870
rect 24872 40769 24900 41074
rect 24952 40928 25004 40934
rect 24952 40870 25004 40876
rect 24858 40760 24914 40769
rect 24858 40695 24914 40704
rect 24676 40384 24728 40390
rect 24676 40326 24728 40332
rect 24768 40384 24820 40390
rect 24768 40326 24820 40332
rect 24400 39840 24452 39846
rect 24400 39782 24452 39788
rect 24308 39364 24360 39370
rect 24308 39306 24360 39312
rect 24320 36689 24348 39306
rect 24306 36680 24362 36689
rect 24306 36615 24362 36624
rect 24216 36100 24268 36106
rect 24216 36042 24268 36048
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 23952 33454 23980 35430
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 24044 33998 24072 34886
rect 24228 34610 24256 36042
rect 24308 35012 24360 35018
rect 24308 34954 24360 34960
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24032 33992 24084 33998
rect 24032 33934 24084 33940
rect 23940 33448 23992 33454
rect 23940 33390 23992 33396
rect 23940 32768 23992 32774
rect 23940 32710 23992 32716
rect 23952 31770 23980 32710
rect 23860 31742 23980 31770
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 27674 23796 28358
rect 23756 27668 23808 27674
rect 23756 27610 23808 27616
rect 23860 27470 23888 31742
rect 23940 31408 23992 31414
rect 23940 31350 23992 31356
rect 23952 30870 23980 31350
rect 23940 30864 23992 30870
rect 23940 30806 23992 30812
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 23952 28762 23980 29038
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 24044 28529 24072 33934
rect 24216 33312 24268 33318
rect 24216 33254 24268 33260
rect 24124 31408 24176 31414
rect 24124 31350 24176 31356
rect 24136 30258 24164 31350
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 24136 28762 24164 29242
rect 24124 28756 24176 28762
rect 24124 28698 24176 28704
rect 24030 28520 24086 28529
rect 24030 28455 24086 28464
rect 24228 28082 24256 33254
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 23676 26382 23704 26930
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23676 25974 23704 26318
rect 23664 25968 23716 25974
rect 23664 25910 23716 25916
rect 24044 24954 24072 27814
rect 24320 27554 24348 34954
rect 24412 32978 24440 39782
rect 24492 39296 24544 39302
rect 24492 39238 24544 39244
rect 24504 38962 24532 39238
rect 24492 38956 24544 38962
rect 24492 38898 24544 38904
rect 24504 34241 24532 38898
rect 24584 38344 24636 38350
rect 24688 38321 24716 40326
rect 24780 40118 24808 40326
rect 24768 40112 24820 40118
rect 24768 40054 24820 40060
rect 24584 38286 24636 38292
rect 24674 38312 24730 38321
rect 24596 36922 24624 38286
rect 24674 38247 24730 38256
rect 24780 37505 24808 40054
rect 24860 40044 24912 40050
rect 24860 39986 24912 39992
rect 24872 39953 24900 39986
rect 24858 39944 24914 39953
rect 24858 39879 24914 39888
rect 24872 39642 24900 39879
rect 24860 39636 24912 39642
rect 24860 39578 24912 39584
rect 24964 38434 24992 40870
rect 25332 39137 25360 41074
rect 25504 39364 25556 39370
rect 25504 39306 25556 39312
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 24872 38406 24992 38434
rect 24766 37496 24822 37505
rect 24766 37431 24822 37440
rect 24584 36916 24636 36922
rect 24584 36858 24636 36864
rect 24768 36780 24820 36786
rect 24768 36722 24820 36728
rect 24584 36576 24636 36582
rect 24584 36518 24636 36524
rect 24596 36174 24624 36518
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24490 34232 24546 34241
rect 24490 34167 24546 34176
rect 24584 33516 24636 33522
rect 24584 33458 24636 33464
rect 24400 32972 24452 32978
rect 24400 32914 24452 32920
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24412 29170 24440 30534
rect 24492 30048 24544 30054
rect 24492 29990 24544 29996
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24400 28484 24452 28490
rect 24400 28426 24452 28432
rect 24136 27526 24348 27554
rect 24136 27334 24164 27526
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24124 27328 24176 27334
rect 24122 27296 24124 27305
rect 24216 27328 24268 27334
rect 24176 27296 24178 27305
rect 24216 27270 24268 27276
rect 24122 27231 24178 27240
rect 24136 26042 24164 27231
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 24124 25424 24176 25430
rect 24124 25366 24176 25372
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23676 23322 23704 24074
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23768 20942 23796 21830
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23676 20505 23704 20810
rect 23754 20632 23810 20641
rect 23754 20567 23810 20576
rect 23662 20496 23718 20505
rect 23662 20431 23718 20440
rect 23768 20346 23796 20567
rect 23860 20534 23888 24006
rect 23952 21162 23980 24686
rect 24044 24070 24072 24890
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 24044 22098 24072 24006
rect 24032 22092 24084 22098
rect 24136 22094 24164 25366
rect 24228 23866 24256 27270
rect 24320 26450 24348 27406
rect 24412 27062 24440 28426
rect 24504 27538 24532 29990
rect 24596 29102 24624 33458
rect 24780 33454 24808 36722
rect 24872 34542 24900 38406
rect 24952 38208 25004 38214
rect 24952 38150 25004 38156
rect 24964 35034 24992 38150
rect 25044 37732 25096 37738
rect 25044 37674 25096 37680
rect 25056 35873 25084 37674
rect 25042 35864 25098 35873
rect 25042 35799 25098 35808
rect 24964 35006 25084 35034
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24860 34400 24912 34406
rect 24860 34342 24912 34348
rect 24872 34202 24900 34342
rect 24860 34196 24912 34202
rect 24860 34138 24912 34144
rect 24768 33448 24820 33454
rect 24768 33390 24820 33396
rect 24780 32586 24808 33390
rect 24688 32558 24808 32586
rect 24688 31482 24716 32558
rect 24860 31952 24912 31958
rect 24860 31894 24912 31900
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24676 31476 24728 31482
rect 24676 31418 24728 31424
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 24780 28422 24808 31622
rect 24872 29714 24900 31894
rect 24964 31278 24992 34886
rect 25056 32842 25084 35006
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24964 29238 24992 30126
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24582 27976 24638 27985
rect 24582 27911 24584 27920
rect 24636 27911 24638 27920
rect 24584 27882 24636 27888
rect 24780 27878 24808 28358
rect 25056 28218 25084 32506
rect 25148 32230 25176 38898
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25228 37256 25280 37262
rect 25228 37198 25280 37204
rect 25240 36378 25268 37198
rect 25332 36854 25360 38694
rect 25412 37120 25464 37126
rect 25412 37062 25464 37068
rect 25320 36848 25372 36854
rect 25320 36790 25372 36796
rect 25228 36372 25280 36378
rect 25228 36314 25280 36320
rect 25228 35080 25280 35086
rect 25228 35022 25280 35028
rect 25240 34202 25268 35022
rect 25320 34536 25372 34542
rect 25320 34478 25372 34484
rect 25228 34196 25280 34202
rect 25228 34138 25280 34144
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 25240 32910 25268 33594
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25136 32224 25188 32230
rect 25136 32166 25188 32172
rect 25044 28212 25096 28218
rect 25044 28154 25096 28160
rect 25148 28014 25176 32166
rect 25332 31890 25360 34478
rect 25424 32366 25452 37062
rect 25412 32360 25464 32366
rect 25412 32302 25464 32308
rect 25412 32020 25464 32026
rect 25412 31962 25464 31968
rect 25320 31884 25372 31890
rect 25320 31826 25372 31832
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25240 30938 25268 31758
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24492 27532 24544 27538
rect 24492 27474 24544 27480
rect 24400 27056 24452 27062
rect 24400 26998 24452 27004
rect 24308 26444 24360 26450
rect 24308 26386 24360 26392
rect 24320 25140 24348 26386
rect 24412 26382 24440 26998
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24504 26058 24532 27474
rect 24952 27328 25004 27334
rect 24950 27296 24952 27305
rect 25004 27296 25006 27305
rect 24950 27231 25006 27240
rect 25240 26994 25268 29446
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25044 26512 25096 26518
rect 25044 26454 25096 26460
rect 24412 26030 24532 26058
rect 24412 25294 24440 26030
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24320 25112 24440 25140
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24136 22066 24348 22094
rect 24032 22034 24084 22040
rect 24044 21350 24072 22034
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 23952 21134 24164 21162
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 23848 20392 23900 20398
rect 23768 20340 23848 20346
rect 23768 20334 23900 20340
rect 23768 20318 23888 20334
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23386 18119 23442 18128
rect 23480 18148 23532 18154
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22848 14600 22876 18022
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22926 17368 22982 17377
rect 22926 17303 22928 17312
rect 22980 17303 22982 17312
rect 22928 17274 22980 17280
rect 23400 17202 23428 18119
rect 23480 18090 23532 18096
rect 23584 17746 23612 18566
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23308 14634 23336 15982
rect 23386 14648 23442 14657
rect 23308 14606 23386 14634
rect 22848 14572 23060 14600
rect 23386 14583 23442 14592
rect 23032 14346 23060 14572
rect 23020 14340 23072 14346
rect 23020 14282 23072 14288
rect 23032 14006 23060 14282
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22848 12782 22876 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22940 12628 22968 13126
rect 23296 12912 23348 12918
rect 23294 12880 23296 12889
rect 23348 12880 23350 12889
rect 23294 12815 23350 12824
rect 22848 12600 22968 12628
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22664 10674 22692 12242
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11354 22784 12174
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22282 3224 22338 3233
rect 22282 3159 22338 3168
rect 22112 2746 22232 2774
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22112 800 22140 2746
rect 22388 2650 22416 8366
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 22190 2408 22246 2417
rect 22190 2343 22246 2352
rect 22204 1834 22232 2343
rect 22192 1828 22244 1834
rect 22192 1770 22244 1776
rect 22296 1601 22324 2586
rect 22282 1592 22338 1601
rect 22282 1527 22338 1536
rect 22480 800 22508 7754
rect 22572 3602 22600 10610
rect 22664 9042 22692 10610
rect 22756 10577 22784 11086
rect 22742 10568 22798 10577
rect 22742 10503 22798 10512
rect 22756 9586 22784 10503
rect 22848 9926 22876 12600
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23492 12374 23520 17070
rect 23676 14618 23704 20198
rect 23754 19680 23810 19689
rect 23754 19615 23810 19624
rect 23768 19514 23796 19615
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23860 17338 23888 20318
rect 23952 19417 23980 20878
rect 24030 19816 24086 19825
rect 24030 19751 24086 19760
rect 23938 19408 23994 19417
rect 23938 19343 23940 19352
rect 23992 19343 23994 19352
rect 23940 19314 23992 19320
rect 24044 19258 24072 19751
rect 23952 19230 24072 19258
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23952 17218 23980 19230
rect 23768 17190 23980 17218
rect 24032 17196 24084 17202
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 23294 11656 23350 11665
rect 23294 11591 23350 11600
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 10742 23336 11591
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23204 10056 23256 10062
rect 23202 10024 23204 10033
rect 23256 10024 23258 10033
rect 23202 9959 23258 9968
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 23308 9602 23336 10678
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23492 10130 23520 10406
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 22744 9580 22796 9586
rect 23308 9574 23428 9602
rect 22744 9522 22796 9528
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22756 7478 22784 8774
rect 22848 7954 22876 8774
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22664 5250 22692 7278
rect 22756 5370 22784 7414
rect 23308 7154 23336 9454
rect 23400 7834 23428 9574
rect 23400 7806 23520 7834
rect 23308 7126 23428 7154
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22664 5222 22784 5250
rect 22652 4616 22704 4622
rect 22650 4584 22652 4593
rect 22704 4584 22706 4593
rect 22650 4519 22706 4528
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22756 2774 22784 5222
rect 22848 4146 22876 5646
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23308 3670 23336 5850
rect 23400 4865 23428 7126
rect 23386 4856 23442 4865
rect 23386 4791 23442 4800
rect 23386 4040 23442 4049
rect 23386 3975 23442 3984
rect 23296 3664 23348 3670
rect 23296 3606 23348 3612
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 22756 2746 22876 2774
rect 22848 800 22876 2746
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 23216 800 23244 2586
rect 23308 1193 23336 3470
rect 23400 3126 23428 3975
rect 23492 3398 23520 7806
rect 23584 5778 23612 11494
rect 23676 11257 23704 14554
rect 23768 13326 23796 17190
rect 24032 17138 24084 17144
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 23952 14074 23980 16050
rect 24044 15162 24072 17138
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23860 12918 23888 13942
rect 23938 13832 23994 13841
rect 23938 13767 23994 13776
rect 23952 13394 23980 13767
rect 24136 13530 24164 21134
rect 24228 18630 24256 21422
rect 24320 19854 24348 22066
rect 24308 19848 24360 19854
rect 24308 19790 24360 19796
rect 24306 18864 24362 18873
rect 24306 18799 24362 18808
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24320 18442 24348 18799
rect 24228 18414 24348 18442
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24228 13410 24256 18414
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 24136 13382 24256 13410
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23938 12880 23994 12889
rect 23860 12782 23888 12854
rect 23938 12815 23994 12824
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23754 11792 23810 11801
rect 23754 11727 23756 11736
rect 23808 11727 23810 11736
rect 23756 11698 23808 11704
rect 23662 11248 23718 11257
rect 23662 11183 23718 11192
rect 23676 11014 23704 11183
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23294 1184 23350 1193
rect 23294 1119 23350 1128
rect 23584 800 23612 4082
rect 23676 3670 23704 9522
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23768 2650 23796 11698
rect 23848 9920 23900 9926
rect 23846 9888 23848 9897
rect 23900 9888 23902 9897
rect 23846 9823 23902 9832
rect 23952 7546 23980 12815
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9722 24072 9862
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23846 7304 23902 7313
rect 23846 7239 23848 7248
rect 23900 7239 23902 7248
rect 23848 7210 23900 7216
rect 24044 5778 24072 7958
rect 24136 7342 24164 13382
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24228 12306 24256 13262
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24320 10062 24348 17206
rect 24412 15026 24440 25112
rect 24596 24206 24624 25638
rect 24950 25256 25006 25265
rect 24950 25191 24952 25200
rect 25004 25191 25006 25200
rect 24952 25162 25004 25168
rect 24766 24440 24822 24449
rect 24766 24375 24822 24384
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24490 23624 24546 23633
rect 24490 23559 24546 23568
rect 24504 23186 24532 23559
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 24504 21706 24532 22034
rect 24582 21992 24638 22001
rect 24582 21927 24638 21936
rect 24596 21894 24624 21927
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24504 21678 24624 21706
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24504 19310 24532 21286
rect 24596 20806 24624 21678
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24688 19514 24716 22918
rect 24780 22574 24808 24375
rect 24858 24032 24914 24041
rect 24858 23967 24914 23976
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24504 14906 24532 19246
rect 24766 18728 24822 18737
rect 24766 18663 24822 18672
rect 24582 17640 24638 17649
rect 24582 17575 24638 17584
rect 24596 17542 24624 17575
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24688 16726 24716 17478
rect 24780 17134 24808 18663
rect 24872 18442 24900 23967
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24964 23769 24992 23802
rect 24950 23760 25006 23769
rect 24950 23695 25006 23704
rect 24950 22808 25006 22817
rect 24950 22743 25006 22752
rect 24964 22642 24992 22743
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 25056 22098 25084 26454
rect 25148 24410 25176 26522
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25332 26194 25360 26386
rect 25424 26382 25452 31962
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25332 26166 25452 26194
rect 25424 25702 25452 26166
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 25240 24886 25268 25638
rect 25228 24880 25280 24886
rect 25280 24840 25360 24868
rect 25228 24822 25280 24828
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 25042 21992 25098 22001
rect 25042 21927 25098 21936
rect 24952 21888 25004 21894
rect 24950 21856 24952 21865
rect 25004 21856 25006 21865
rect 24950 21791 25006 21800
rect 24952 21072 25004 21078
rect 24952 21014 25004 21020
rect 24964 20618 24992 21014
rect 25056 21010 25084 21927
rect 25148 21146 25176 23122
rect 25240 22098 25268 24550
rect 25332 24138 25360 24840
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25332 23798 25360 24074
rect 25424 23866 25452 25638
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25332 22438 25360 23734
rect 25410 22536 25466 22545
rect 25410 22471 25466 22480
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25044 21004 25096 21010
rect 25044 20946 25096 20952
rect 24964 20590 25084 20618
rect 24950 20360 25006 20369
rect 24950 20295 25006 20304
rect 24964 19922 24992 20295
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 24872 18414 24992 18442
rect 24858 17912 24914 17921
rect 24858 17847 24914 17856
rect 24872 17746 24900 17847
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24674 15192 24730 15201
rect 24674 15127 24730 15136
rect 24688 15026 24716 15127
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24504 14878 24716 14906
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24504 13258 24532 13806
rect 24584 13320 24636 13326
rect 24582 13288 24584 13297
rect 24636 13288 24638 13297
rect 24492 13252 24544 13258
rect 24582 13223 24638 13232
rect 24492 13194 24544 13200
rect 24504 12900 24532 13194
rect 24584 12912 24636 12918
rect 24504 12872 24584 12900
rect 24584 12854 24636 12860
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 12434 24532 12718
rect 24412 12406 24532 12434
rect 24412 10674 24440 12406
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24308 10056 24360 10062
rect 24308 9998 24360 10004
rect 24412 7834 24440 10610
rect 24320 7806 24440 7834
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 23938 5264 23994 5273
rect 23938 5199 23940 5208
rect 23992 5199 23994 5208
rect 23940 5170 23992 5176
rect 24320 4282 24348 7806
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23860 3738 23888 4082
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23846 3632 23902 3641
rect 23846 3567 23902 3576
rect 23860 3058 23888 3567
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23952 800 23980 4082
rect 24214 3768 24270 3777
rect 24214 3703 24216 3712
rect 24268 3703 24270 3712
rect 24216 3674 24268 3680
rect 24320 3534 24348 4218
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 2582 24256 3402
rect 24216 2576 24268 2582
rect 24216 2518 24268 2524
rect 24412 1358 24440 7686
rect 24504 5710 24532 10950
rect 24688 8974 24716 14878
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24766 13016 24822 13025
rect 24766 12951 24822 12960
rect 24780 11694 24808 12951
rect 24872 12850 24900 13670
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24858 12200 24914 12209
rect 24858 12135 24914 12144
rect 24872 11830 24900 12135
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24872 11082 24900 11319
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24766 10568 24822 10577
rect 24766 10503 24822 10512
rect 24780 9518 24808 10503
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24858 8936 24914 8945
rect 24858 8871 24914 8880
rect 24872 8430 24900 8871
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24858 8120 24914 8129
rect 24858 8055 24914 8064
rect 24872 7954 24900 8055
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24766 7304 24822 7313
rect 24766 7239 24822 7248
rect 24674 6896 24730 6905
rect 24674 6831 24730 6840
rect 24688 6798 24716 6831
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24780 6254 24808 7239
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24582 5672 24638 5681
rect 24582 5607 24638 5616
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24596 5574 24624 5607
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24780 5166 24808 5607
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24504 2650 24532 3470
rect 24596 2650 24624 4558
rect 24964 4146 24992 18414
rect 25056 17746 25084 20590
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 25148 19718 25176 20470
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 25136 19304 25188 19310
rect 25134 19272 25136 19281
rect 25188 19272 25190 19281
rect 25134 19207 25190 19216
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25148 17202 25176 18022
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25134 17096 25190 17105
rect 25134 17031 25190 17040
rect 25044 16516 25096 16522
rect 25044 16458 25096 16464
rect 25056 16289 25084 16458
rect 25042 16280 25098 16289
rect 25042 16215 25098 16224
rect 25148 16182 25176 17031
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 25240 15502 25268 22034
rect 25228 15496 25280 15502
rect 25042 15464 25098 15473
rect 25228 15438 25280 15444
rect 25042 15399 25044 15408
rect 25096 15399 25098 15408
rect 25044 15370 25096 15376
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 25056 12238 25084 14214
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 25056 10742 25084 10950
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 25148 10690 25176 14350
rect 25240 13938 25268 15302
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 25240 10826 25268 13738
rect 25332 12442 25360 22170
rect 25424 13802 25452 22471
rect 25516 21350 25544 39306
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 25596 33856 25648 33862
rect 25596 33798 25648 33804
rect 25608 23118 25636 33798
rect 25700 25498 25728 33934
rect 25792 29306 25820 47398
rect 26148 40384 26200 40390
rect 26148 40326 26200 40332
rect 25872 35624 25924 35630
rect 25872 35566 25924 35572
rect 25884 33658 25912 35566
rect 25872 33652 25924 33658
rect 25872 33594 25924 33600
rect 25780 29300 25832 29306
rect 25780 29242 25832 29248
rect 25884 28642 25912 33594
rect 26160 31142 26188 40326
rect 26148 31136 26200 31142
rect 26148 31078 26200 31084
rect 25964 30864 26016 30870
rect 25964 30806 26016 30812
rect 25792 28614 25912 28642
rect 25792 28490 25820 28614
rect 25976 28506 26004 30806
rect 25780 28484 25832 28490
rect 25780 28426 25832 28432
rect 25884 28478 26004 28506
rect 25780 26308 25832 26314
rect 25780 26250 25832 26256
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25688 23656 25740 23662
rect 25688 23598 25740 23604
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25608 21622 25636 22374
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25516 20602 25544 21082
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25516 19514 25544 20538
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25412 13796 25464 13802
rect 25412 13738 25464 13744
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25240 10798 25360 10826
rect 25148 10662 25268 10690
rect 25134 9752 25190 9761
rect 25134 9687 25190 9696
rect 25148 8566 25176 9687
rect 25240 9178 25268 10662
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25332 7274 25360 10798
rect 25320 7268 25372 7274
rect 25320 7210 25372 7216
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 25056 6497 25084 6666
rect 25042 6488 25098 6497
rect 25042 6423 25098 6432
rect 25332 5778 25360 7210
rect 25516 6866 25544 18566
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25608 8090 25636 18158
rect 25700 10266 25728 23598
rect 25792 23050 25820 26250
rect 25780 23044 25832 23050
rect 25780 22986 25832 22992
rect 25884 22094 25912 28478
rect 25964 26920 26016 26926
rect 25964 26862 26016 26868
rect 25792 22066 25912 22094
rect 25792 14074 25820 22066
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25884 15337 25912 21286
rect 25976 16590 26004 26862
rect 26148 23044 26200 23050
rect 26148 22986 26200 22992
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26068 18970 26096 22442
rect 26160 19310 26188 22986
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 25870 15328 25926 15337
rect 25870 15263 25926 15272
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24596 1562 24624 2382
rect 24584 1556 24636 1562
rect 24584 1498 24636 1504
rect 24400 1352 24452 1358
rect 24400 1294 24452 1300
rect 24228 870 24348 898
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24228 134 24256 870
rect 24320 800 24348 870
rect 24216 128 24268 134
rect 24216 70 24268 76
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24964 785 24992 3878
rect 24950 776 25006 785
rect 24950 711 25006 720
rect 25042 0 25098 800
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 4342 29008 4398 29064
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 3974 19896 4030 19952
rect 5538 27376 5594 27432
rect 7194 23604 7196 23624
rect 7196 23604 7248 23624
rect 7248 23604 7250 23624
rect 7194 23568 7250 23604
rect 4618 19796 4620 19816
rect 4620 19796 4672 19816
rect 4672 19796 4674 19816
rect 4618 19760 4674 19796
rect 1306 17720 1362 17776
rect 1766 15544 1822 15600
rect 2042 15308 2044 15328
rect 2044 15308 2096 15328
rect 2096 15308 2098 15328
rect 2042 15272 2098 15308
rect 1858 13912 1914 13968
rect 1766 12708 1822 12744
rect 1766 12688 1768 12708
rect 1768 12688 1820 12708
rect 1820 12688 1822 12708
rect 1490 7656 1546 7712
rect 1306 5480 1362 5536
rect 1858 9460 1860 9480
rect 1860 9460 1912 9480
rect 1912 9460 1914 9480
rect 1858 9424 1914 9460
rect 2042 14184 2098 14240
rect 2134 12280 2190 12336
rect 2134 12180 2136 12200
rect 2136 12180 2188 12200
rect 2188 12180 2190 12200
rect 2134 12144 2190 12180
rect 2042 10920 2098 10976
rect 2042 9696 2098 9752
rect 1950 8336 2006 8392
rect 1674 4528 1730 4584
rect 1674 3984 1730 4040
rect 1858 3168 1914 3224
rect 2410 7928 2466 7984
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 4066 18672 4122 18728
rect 5170 21392 5226 21448
rect 5078 19352 5134 19408
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 3422 15680 3478 15736
rect 2594 13776 2650 13832
rect 2686 10104 2742 10160
rect 2686 9832 2742 9888
rect 2686 8356 2742 8392
rect 2686 8336 2688 8356
rect 2688 8336 2740 8356
rect 2740 8336 2742 8356
rect 3238 14864 3294 14920
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 3238 11076 3294 11112
rect 3238 11056 3240 11076
rect 3240 11056 3292 11076
rect 3292 11056 3294 11076
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3238 9988 3294 10024
rect 3238 9968 3240 9988
rect 3240 9968 3292 9988
rect 3292 9968 3294 9988
rect 3238 9596 3240 9616
rect 3240 9596 3292 9616
rect 3292 9596 3294 9616
rect 3238 9560 3294 9596
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3238 4664 3294 4720
rect 2870 4120 2926 4176
rect 2870 3984 2926 4040
rect 3422 13640 3478 13696
rect 4526 17856 4582 17912
rect 4066 15952 4122 16008
rect 3606 12416 3662 12472
rect 3606 10548 3608 10568
rect 3608 10548 3660 10568
rect 3660 10548 3662 10568
rect 3606 10512 3662 10548
rect 3606 10376 3662 10432
rect 3422 9016 3478 9072
rect 3514 8064 3570 8120
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2318 1672 2374 1728
rect 2686 3304 2742 3360
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3790 14728 3846 14784
rect 3790 13912 3846 13968
rect 3790 12588 3792 12608
rect 3792 12588 3844 12608
rect 3844 12588 3846 12608
rect 3790 12552 3846 12588
rect 4066 13912 4122 13968
rect 4250 15428 4306 15464
rect 4250 15408 4252 15428
rect 4252 15408 4304 15428
rect 4304 15408 4306 15428
rect 4434 15816 4490 15872
rect 4250 13368 4306 13424
rect 4066 12300 4122 12336
rect 4066 12280 4068 12300
rect 4068 12280 4120 12300
rect 4120 12280 4122 12300
rect 3974 11756 4030 11792
rect 3974 11736 3976 11756
rect 3976 11736 4028 11756
rect 4028 11736 4030 11756
rect 3974 8880 4030 8936
rect 4066 8744 4122 8800
rect 4250 10240 4306 10296
rect 3974 8064 4030 8120
rect 4066 6740 4068 6760
rect 4068 6740 4120 6760
rect 4120 6740 4122 6760
rect 4066 6704 4122 6740
rect 4158 5636 4214 5672
rect 4158 5616 4160 5636
rect 4160 5616 4212 5636
rect 4212 5616 4214 5636
rect 3882 3052 3938 3088
rect 3882 3032 3884 3052
rect 3884 3032 3936 3052
rect 3936 3032 3938 3052
rect 4066 4256 4122 4312
rect 4434 7928 4490 7984
rect 4342 7404 4398 7440
rect 4342 7384 4344 7404
rect 4344 7384 4396 7404
rect 4396 7384 4398 7404
rect 4342 6196 4344 6216
rect 4344 6196 4396 6216
rect 4396 6196 4398 6216
rect 4342 6160 4398 6196
rect 4710 18164 4712 18184
rect 4712 18164 4764 18184
rect 4764 18164 4766 18184
rect 4710 18128 4766 18164
rect 4894 17176 4950 17232
rect 4710 17040 4766 17096
rect 4986 16088 5042 16144
rect 5078 15408 5134 15464
rect 5354 20032 5410 20088
rect 6274 23160 6330 23216
rect 6182 19216 6238 19272
rect 5722 18808 5778 18864
rect 5262 14340 5318 14376
rect 5262 14320 5264 14340
rect 5264 14320 5316 14340
rect 5316 14320 5318 14340
rect 6090 17584 6146 17640
rect 5170 13252 5226 13288
rect 5170 13232 5172 13252
rect 5172 13232 5224 13252
rect 5224 13232 5226 13252
rect 5078 12844 5134 12880
rect 5078 12824 5080 12844
rect 5080 12824 5132 12844
rect 5132 12824 5134 12844
rect 4986 9868 4988 9888
rect 4988 9868 5040 9888
rect 5040 9868 5042 9888
rect 4986 9832 5042 9868
rect 4986 8744 5042 8800
rect 4986 8200 5042 8256
rect 4894 7656 4950 7712
rect 4894 7148 4896 7168
rect 4896 7148 4948 7168
rect 4948 7148 4950 7168
rect 4894 7112 4950 7148
rect 4894 6976 4950 7032
rect 4618 3712 4674 3768
rect 5538 12688 5594 12744
rect 5630 12552 5686 12608
rect 5446 8880 5502 8936
rect 5262 8472 5318 8528
rect 5078 6296 5134 6352
rect 5170 5888 5226 5944
rect 5446 2508 5502 2544
rect 5446 2488 5448 2508
rect 5448 2488 5500 2508
rect 5500 2488 5502 2508
rect 5722 5344 5778 5400
rect 5630 4800 5686 4856
rect 6550 21936 6606 21992
rect 6734 20440 6790 20496
rect 6458 16632 6514 16688
rect 5998 11636 6000 11656
rect 6000 11636 6052 11656
rect 6052 11636 6054 11656
rect 5998 11600 6054 11636
rect 5906 8608 5962 8664
rect 5906 7248 5962 7304
rect 5906 3984 5962 4040
rect 7378 20168 7434 20224
rect 7378 16768 7434 16824
rect 6274 14456 6330 14512
rect 6182 12552 6238 12608
rect 6090 3984 6146 4040
rect 6550 14884 6606 14920
rect 6550 14864 6552 14884
rect 6552 14864 6604 14884
rect 6604 14864 6606 14884
rect 6550 14592 6606 14648
rect 7194 15000 7250 15056
rect 6918 13776 6974 13832
rect 6642 12588 6644 12608
rect 6644 12588 6696 12608
rect 6696 12588 6698 12608
rect 6642 12552 6698 12588
rect 6918 11464 6974 11520
rect 6458 6976 6514 7032
rect 6642 10104 6698 10160
rect 6826 8880 6882 8936
rect 6826 7384 6882 7440
rect 6642 6976 6698 7032
rect 6182 2932 6184 2952
rect 6184 2932 6236 2952
rect 6236 2932 6238 2952
rect 6182 2896 6238 2932
rect 6366 2352 6422 2408
rect 6642 3576 6698 3632
rect 7562 15136 7618 15192
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 8942 24656 8998 24712
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8114 20476 8116 20496
rect 8116 20476 8168 20496
rect 8168 20476 8170 20496
rect 8114 20440 8170 20476
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8390 20304 8446 20360
rect 8666 20032 8722 20088
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 9126 22072 9182 22128
rect 8666 19760 8722 19816
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7930 16496 7986 16552
rect 8298 16668 8300 16688
rect 8300 16668 8352 16688
rect 8352 16668 8354 16688
rect 8298 16632 8354 16668
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8482 16396 8484 16416
rect 8484 16396 8536 16416
rect 8536 16396 8538 16416
rect 8482 16360 8538 16396
rect 7930 15408 7986 15464
rect 8114 15408 8170 15464
rect 8390 15544 8446 15600
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7930 15000 7986 15056
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7562 12416 7618 12472
rect 7010 10240 7066 10296
rect 7470 11192 7526 11248
rect 7286 10684 7288 10704
rect 7288 10684 7340 10704
rect 7340 10684 7342 10704
rect 7286 10648 7342 10684
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 8390 15272 8446 15328
rect 8298 11328 8354 11384
rect 9034 19488 9090 19544
rect 10138 29416 10194 29472
rect 9310 27276 9312 27296
rect 9312 27276 9364 27296
rect 9364 27276 9366 27296
rect 9310 27240 9366 27276
rect 9218 17992 9274 18048
rect 9678 18264 9734 18320
rect 9034 16224 9090 16280
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7010 7112 7066 7168
rect 7286 7792 7342 7848
rect 7102 6840 7158 6896
rect 6826 1400 6882 1456
rect 7286 5616 7342 5672
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 8758 12416 8814 12472
rect 8482 10648 8538 10704
rect 8206 9288 8262 9344
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 8482 9152 8538 9208
rect 7930 8064 7986 8120
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7654 5772 7710 5808
rect 7654 5752 7656 5772
rect 7656 5752 7708 5772
rect 7708 5752 7710 5772
rect 7562 5480 7618 5536
rect 7470 3440 7526 3496
rect 7654 5364 7710 5400
rect 7654 5344 7656 5364
rect 7656 5344 7708 5364
rect 7708 5344 7710 5364
rect 7654 5208 7710 5264
rect 7930 5616 7986 5672
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 8298 4664 8354 4720
rect 8574 7520 8630 7576
rect 8574 6840 8630 6896
rect 8574 6568 8630 6624
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 8482 4392 8538 4448
rect 8390 4256 8446 4312
rect 7654 3304 7710 3360
rect 7654 3168 7710 3224
rect 7930 3576 7986 3632
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 8298 2796 8300 2816
rect 8300 2796 8352 2816
rect 8352 2796 8354 2816
rect 8298 2760 8354 2796
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 7930 1300 7932 1320
rect 7932 1300 7984 1320
rect 7984 1300 7986 1320
rect 7930 1264 7986 1300
rect 8390 2624 8446 2680
rect 8390 2080 8446 2136
rect 9954 18400 10010 18456
rect 9770 17720 9826 17776
rect 9954 17448 10010 17504
rect 10322 26460 10324 26480
rect 10324 26460 10376 26480
rect 10376 26460 10378 26480
rect 10322 26424 10378 26460
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 10966 27920 11022 27976
rect 10598 26016 10654 26072
rect 10138 17720 10194 17776
rect 9770 16632 9826 16688
rect 10138 16904 10194 16960
rect 9954 16244 10010 16280
rect 9954 16224 9956 16244
rect 9956 16224 10008 16244
rect 10008 16224 10010 16244
rect 9954 13504 10010 13560
rect 9770 12960 9826 13016
rect 10138 12416 10194 12472
rect 9678 12008 9734 12064
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 11242 15816 11298 15872
rect 10874 15136 10930 15192
rect 10874 14068 10930 14104
rect 10874 14048 10876 14068
rect 10876 14048 10928 14068
rect 10928 14048 10930 14068
rect 10506 11872 10562 11928
rect 10322 11464 10378 11520
rect 8850 9036 8906 9072
rect 8850 9016 8852 9036
rect 8852 9016 8904 9036
rect 8904 9016 8906 9036
rect 8942 8064 8998 8120
rect 8758 5616 8814 5672
rect 8850 4256 8906 4312
rect 9586 9868 9588 9888
rect 9588 9868 9640 9888
rect 9640 9868 9642 9888
rect 9586 9832 9642 9868
rect 10414 9696 10470 9752
rect 10598 10784 10654 10840
rect 11518 16904 11574 16960
rect 11334 14728 11390 14784
rect 11242 14184 11298 14240
rect 10230 8608 10286 8664
rect 9586 7828 9588 7848
rect 9588 7828 9640 7848
rect 9640 7828 9642 7848
rect 9586 7792 9642 7828
rect 9126 4936 9182 4992
rect 8758 3304 8814 3360
rect 8942 2896 8998 2952
rect 9310 5072 9366 5128
rect 9678 4156 9680 4176
rect 9680 4156 9732 4176
rect 9732 4156 9734 4176
rect 9678 4120 9734 4156
rect 11242 7520 11298 7576
rect 11978 20576 12034 20632
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12714 29688 12770 29744
rect 13542 29552 13598 29608
rect 12990 29452 12992 29472
rect 12992 29452 13044 29472
rect 13044 29452 13046 29472
rect 12990 29416 13046 29452
rect 13818 29280 13874 29336
rect 13726 29144 13782 29200
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 13726 26696 13782 26752
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12622 24148 12624 24168
rect 12624 24148 12676 24168
rect 12676 24148 12678 24168
rect 12622 24112 12678 24148
rect 13266 23840 13322 23896
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13450 24012 13452 24032
rect 13452 24012 13504 24032
rect 13504 24012 13506 24032
rect 13450 23976 13506 24012
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12438 20168 12494 20224
rect 11794 17992 11850 18048
rect 11978 17992 12034 18048
rect 11886 16904 11942 16960
rect 11702 12960 11758 13016
rect 12254 16360 12310 16416
rect 12070 13252 12126 13288
rect 12070 13232 12072 13252
rect 12072 13232 12124 13252
rect 12124 13232 12126 13252
rect 11702 12416 11758 12472
rect 11610 12280 11666 12336
rect 11426 10376 11482 10432
rect 11610 10240 11666 10296
rect 11334 6840 11390 6896
rect 10966 5208 11022 5264
rect 11058 3712 11114 3768
rect 11978 11872 12034 11928
rect 11794 10412 11796 10432
rect 11796 10412 11848 10432
rect 11848 10412 11850 10432
rect 11794 10376 11850 10412
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 14002 23740 14004 23760
rect 14004 23740 14056 23760
rect 14056 23740 14058 23760
rect 14002 23704 14058 23740
rect 13634 21120 13690 21176
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12162 12416 12218 12472
rect 12346 12960 12402 13016
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 14278 23432 14334 23488
rect 14462 27240 14518 27296
rect 14462 25472 14518 25528
rect 14186 20748 14188 20768
rect 14188 20748 14240 20768
rect 14240 20748 14242 20768
rect 14186 20712 14242 20748
rect 14738 27276 14740 27296
rect 14740 27276 14792 27296
rect 14792 27276 14794 27296
rect 14738 27240 14794 27276
rect 14646 23976 14702 24032
rect 15106 29300 15162 29336
rect 15106 29280 15108 29300
rect 15108 29280 15160 29300
rect 15160 29280 15162 29300
rect 15290 29708 15346 29744
rect 15290 29688 15292 29708
rect 15292 29688 15344 29708
rect 15344 29688 15346 29708
rect 15290 28600 15346 28656
rect 15658 28872 15714 28928
rect 14830 24112 14886 24168
rect 15106 23432 15162 23488
rect 14370 20032 14426 20088
rect 16026 29416 16082 29472
rect 15934 28620 15990 28656
rect 15934 28600 15936 28620
rect 15936 28600 15988 28620
rect 15988 28600 15990 28620
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 22374 55392 22430 55448
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17038 35808 17094 35864
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17314 34448 17370 34504
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 16302 27276 16304 27296
rect 16304 27276 16356 27296
rect 16356 27276 16358 27296
rect 16302 27240 16358 27276
rect 14554 19488 14610 19544
rect 14186 18028 14188 18048
rect 14188 18028 14240 18048
rect 14240 18028 14242 18048
rect 14186 17992 14242 18028
rect 14002 16224 14058 16280
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13358 13676 13360 13696
rect 13360 13676 13412 13696
rect 13412 13676 13414 13696
rect 13358 13640 13414 13676
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13726 12552 13782 12608
rect 13634 12316 13636 12336
rect 13636 12316 13688 12336
rect 13688 12316 13690 12336
rect 13634 12280 13690 12316
rect 12714 11464 12770 11520
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13634 11328 13690 11384
rect 12714 10376 12770 10432
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13174 9696 13230 9752
rect 12254 8608 12310 8664
rect 12346 6840 12402 6896
rect 12162 6024 12218 6080
rect 11978 5888 12034 5944
rect 11886 5480 11942 5536
rect 11794 4528 11850 4584
rect 12346 5888 12402 5944
rect 12346 4800 12402 4856
rect 12346 4528 12402 4584
rect 12622 6860 12678 6896
rect 12622 6840 12624 6860
rect 12624 6840 12676 6860
rect 12676 6840 12678 6860
rect 12530 6432 12586 6488
rect 12622 6024 12678 6080
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13266 8472 13322 8528
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12806 8064 12862 8120
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 14830 20576 14886 20632
rect 13818 9696 13874 9752
rect 13542 8064 13598 8120
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13542 6432 13598 6488
rect 13542 5908 13598 5944
rect 13542 5888 13544 5908
rect 13544 5888 13596 5908
rect 13596 5888 13598 5908
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12622 3984 12678 4040
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12530 1672 12586 1728
rect 13450 3848 13506 3904
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 13910 4936 13966 4992
rect 13542 1944 13598 2000
rect 14830 15136 14886 15192
rect 15290 19080 15346 19136
rect 15106 18536 15162 18592
rect 15474 17312 15530 17368
rect 15290 15972 15346 16008
rect 15290 15952 15292 15972
rect 15292 15952 15344 15972
rect 15344 15952 15346 15972
rect 15198 15544 15254 15600
rect 15198 13776 15254 13832
rect 14186 9288 14242 9344
rect 14462 10240 14518 10296
rect 14370 9288 14426 9344
rect 14462 8064 14518 8120
rect 14278 7692 14280 7712
rect 14280 7692 14332 7712
rect 14332 7692 14334 7712
rect 14278 7656 14334 7692
rect 14922 12008 14978 12064
rect 15566 15544 15622 15600
rect 15474 13504 15530 13560
rect 15474 12960 15530 13016
rect 14922 10240 14978 10296
rect 14278 4800 14334 4856
rect 14738 6568 14794 6624
rect 14922 6840 14978 6896
rect 14922 6568 14978 6624
rect 14738 5480 14794 5536
rect 14922 5344 14978 5400
rect 14462 3712 14518 3768
rect 14094 2488 14150 2544
rect 15566 12552 15622 12608
rect 16118 25336 16174 25392
rect 17130 26424 17186 26480
rect 15750 17876 15806 17912
rect 15750 17856 15752 17876
rect 15752 17856 15804 17876
rect 15804 17856 15806 17876
rect 16486 23704 16542 23760
rect 16394 23568 16450 23624
rect 16394 22616 16450 22672
rect 16394 22516 16396 22536
rect 16396 22516 16448 22536
rect 16448 22516 16450 22536
rect 16394 22480 16450 22516
rect 16394 21392 16450 21448
rect 16118 16632 16174 16688
rect 15934 15272 15990 15328
rect 17498 28872 17554 28928
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 18602 30776 18658 30832
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17130 21392 17186 21448
rect 17038 19352 17094 19408
rect 16302 17992 16358 18048
rect 16394 17448 16450 17504
rect 16394 16632 16450 16688
rect 16670 16088 16726 16144
rect 15842 13504 15898 13560
rect 16118 13640 16174 13696
rect 15474 6604 15476 6624
rect 15476 6604 15528 6624
rect 15528 6604 15530 6624
rect 15474 6568 15530 6604
rect 15474 6432 15530 6488
rect 16118 12960 16174 13016
rect 16394 14184 16450 14240
rect 16486 14048 16542 14104
rect 16486 13776 16542 13832
rect 16394 12416 16450 12472
rect 16486 12144 16542 12200
rect 16302 10920 16358 10976
rect 16578 12008 16634 12064
rect 16578 11192 16634 11248
rect 16394 9832 16450 9888
rect 16026 9288 16082 9344
rect 15750 8472 15806 8528
rect 15566 5752 15622 5808
rect 15106 3304 15162 3360
rect 15290 1400 15346 1456
rect 15934 8336 15990 8392
rect 15934 6860 15990 6896
rect 15934 6840 15936 6860
rect 15936 6840 15988 6860
rect 15988 6840 15990 6860
rect 15842 6568 15898 6624
rect 15842 6432 15898 6488
rect 16854 16088 16910 16144
rect 17498 20576 17554 20632
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 18050 25764 18106 25800
rect 18050 25744 18052 25764
rect 18052 25744 18104 25764
rect 18104 25744 18106 25764
rect 18694 29552 18750 29608
rect 18786 27512 18842 27568
rect 18694 26424 18750 26480
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 18510 24676 18566 24712
rect 18510 24656 18512 24676
rect 18512 24656 18564 24676
rect 18564 24656 18566 24676
rect 17682 20576 17738 20632
rect 17590 19760 17646 19816
rect 16854 14184 16910 14240
rect 16946 9596 16948 9616
rect 16948 9596 17000 9616
rect 17000 9596 17002 9616
rect 16946 9560 17002 9596
rect 17222 11736 17278 11792
rect 17498 16632 17554 16688
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18326 20052 18382 20088
rect 18326 20032 18328 20052
rect 18328 20032 18380 20052
rect 18380 20032 18382 20052
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 19062 29144 19118 29200
rect 18970 26324 18972 26344
rect 18972 26324 19024 26344
rect 19024 26324 19026 26344
rect 18970 26288 19026 26324
rect 18786 22480 18842 22536
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17866 17176 17922 17232
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18510 15952 18566 16008
rect 18510 15408 18566 15464
rect 17498 12280 17554 12336
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17774 13640 17830 13696
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 19522 23432 19578 23488
rect 18970 20440 19026 20496
rect 19338 21800 19394 21856
rect 19338 20984 19394 21040
rect 19430 20848 19486 20904
rect 18786 17856 18842 17912
rect 18694 16496 18750 16552
rect 19062 17740 19118 17776
rect 19062 17720 19064 17740
rect 19064 17720 19116 17740
rect 19116 17720 19118 17740
rect 18326 12416 18382 12472
rect 17682 12008 17738 12064
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17866 11348 17922 11384
rect 17866 11328 17868 11348
rect 17868 11328 17920 11348
rect 17920 11328 17922 11348
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17866 10104 17922 10160
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 16486 7520 16542 7576
rect 16486 6840 16542 6896
rect 16762 6432 16818 6488
rect 16762 6024 16818 6080
rect 16670 5344 16726 5400
rect 17130 5888 17186 5944
rect 17498 7928 17554 7984
rect 17590 6976 17646 7032
rect 17590 6840 17646 6896
rect 17038 1264 17094 1320
rect 17038 856 17094 912
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18234 6840 18290 6896
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18142 5888 18198 5944
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18510 8336 18566 8392
rect 18694 11056 18750 11112
rect 18694 9016 18750 9072
rect 18694 8336 18750 8392
rect 19062 15680 19118 15736
rect 18970 11212 19026 11248
rect 18970 11192 18972 11212
rect 18972 11192 19024 11212
rect 19024 11192 19026 11212
rect 19614 21800 19670 21856
rect 24122 56208 24178 56264
rect 22834 54576 22890 54632
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 23386 53760 23442 53816
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 21822 32544 21878 32600
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 24582 52944 24638 53000
rect 24950 52128 25006 52184
rect 24950 51332 25006 51368
rect 24950 51312 24952 51332
rect 24952 51312 25004 51332
rect 25004 51312 25006 51332
rect 24950 50496 25006 50552
rect 24766 47640 24822 47696
rect 24858 46960 24914 47016
rect 25502 49680 25558 49736
rect 25134 48864 25190 48920
rect 25134 48084 25136 48104
rect 25136 48084 25188 48104
rect 25188 48084 25190 48104
rect 25134 48048 25190 48084
rect 25226 47504 25282 47560
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 25318 45600 25374 45656
rect 25318 44820 25320 44840
rect 25320 44820 25372 44840
rect 25372 44820 25374 44840
rect 25318 44784 25374 44820
rect 24766 43968 24822 44024
rect 25502 43152 25558 43208
rect 25226 42608 25282 42664
rect 25134 42336 25190 42392
rect 24858 41520 24914 41576
rect 25134 41540 25190 41576
rect 25134 41520 25136 41540
rect 25136 41520 25188 41540
rect 25188 41520 25190 41540
rect 23478 40024 23534 40080
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22742 34992 22798 35048
rect 22098 33360 22154 33416
rect 20718 25336 20774 25392
rect 20810 24928 20866 24984
rect 20442 23976 20498 24032
rect 22098 31728 22154 31784
rect 22098 31184 22154 31240
rect 20994 23432 21050 23488
rect 20810 20748 20812 20768
rect 20812 20748 20864 20768
rect 20864 20748 20866 20768
rect 19522 15272 19578 15328
rect 19338 13524 19394 13560
rect 19338 13504 19340 13524
rect 19340 13504 19392 13524
rect 19392 13504 19394 13524
rect 19522 13096 19578 13152
rect 19338 11348 19394 11384
rect 19338 11328 19340 11348
rect 19340 11328 19392 11348
rect 19392 11328 19394 11348
rect 19154 10648 19210 10704
rect 17774 3576 17830 3632
rect 17406 1128 17462 1184
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18050 3984 18106 4040
rect 18418 5072 18474 5128
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18510 2896 18566 2952
rect 17866 2352 17922 2408
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 16302 448 16358 504
rect 18694 856 18750 912
rect 18878 2896 18934 2952
rect 19338 7112 19394 7168
rect 19338 5888 19394 5944
rect 19246 4936 19302 4992
rect 19154 2896 19210 2952
rect 19430 4120 19486 4176
rect 19798 14728 19854 14784
rect 19706 11464 19762 11520
rect 19982 9424 20038 9480
rect 19614 7928 19670 7984
rect 20810 20712 20866 20748
rect 20810 19896 20866 19952
rect 20718 19760 20774 19816
rect 20626 19624 20682 19680
rect 20350 15000 20406 15056
rect 20442 13932 20498 13968
rect 20442 13912 20444 13932
rect 20444 13912 20496 13932
rect 20496 13912 20498 13932
rect 20810 18672 20866 18728
rect 21270 20848 21326 20904
rect 20626 13388 20682 13424
rect 20626 13368 20628 13388
rect 20628 13368 20680 13388
rect 20680 13368 20682 13388
rect 20718 13232 20774 13288
rect 20718 12588 20720 12608
rect 20720 12588 20772 12608
rect 20772 12588 20774 12608
rect 20718 12552 20774 12588
rect 20902 15272 20958 15328
rect 22006 29028 22062 29064
rect 22006 29008 22008 29028
rect 22008 29008 22060 29028
rect 22060 29008 22062 29028
rect 21822 24928 21878 24984
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22282 26832 22338 26888
rect 22466 26696 22522 26752
rect 22374 26016 22430 26072
rect 22006 23568 22062 23624
rect 22098 23160 22154 23216
rect 21914 22072 21970 22128
rect 21914 21800 21970 21856
rect 21822 20884 21824 20904
rect 21824 20884 21876 20904
rect 21876 20884 21878 20904
rect 21822 20848 21878 20884
rect 22006 21664 22062 21720
rect 22190 21564 22192 21584
rect 22192 21564 22244 21584
rect 22244 21564 22246 21584
rect 22190 21528 22246 21564
rect 22006 20324 22062 20360
rect 22006 20304 22008 20324
rect 22008 20304 22060 20324
rect 22060 20304 22062 20324
rect 22466 21428 22468 21448
rect 22468 21428 22520 21448
rect 22520 21428 22522 21448
rect 22466 21392 22522 21428
rect 21914 18264 21970 18320
rect 21638 14864 21694 14920
rect 21270 14320 21326 14376
rect 20994 12416 21050 12472
rect 20166 11212 20222 11248
rect 20166 11192 20168 11212
rect 20168 11192 20220 11212
rect 20220 11192 20222 11212
rect 20258 9832 20314 9888
rect 19890 7112 19946 7168
rect 19614 6060 19616 6080
rect 19616 6060 19668 6080
rect 19668 6060 19670 6080
rect 19614 6024 19670 6060
rect 19706 5888 19762 5944
rect 19706 4020 19708 4040
rect 19708 4020 19760 4040
rect 19760 4020 19762 4040
rect 19706 3984 19762 4020
rect 20074 6724 20130 6760
rect 20074 6704 20076 6724
rect 20076 6704 20128 6724
rect 20128 6704 20130 6724
rect 19982 5072 20038 5128
rect 19890 3848 19946 3904
rect 20258 7948 20314 7984
rect 20258 7928 20260 7948
rect 20260 7928 20312 7948
rect 20312 7928 20314 7948
rect 20626 8472 20682 8528
rect 20718 7792 20774 7848
rect 20810 6160 20866 6216
rect 20718 4664 20774 4720
rect 21086 9560 21142 9616
rect 20626 3984 20682 4040
rect 20350 1944 20406 2000
rect 21454 12688 21510 12744
rect 21730 14592 21786 14648
rect 22006 14340 22062 14376
rect 22006 14320 22008 14340
rect 22008 14320 22060 14340
rect 22060 14320 22062 14340
rect 22098 12960 22154 13016
rect 21638 11076 21694 11112
rect 21638 11056 21640 11076
rect 21640 11056 21692 11076
rect 21692 11056 21694 11076
rect 21178 4800 21234 4856
rect 20810 992 20866 1048
rect 21730 9560 21786 9616
rect 21638 1808 21694 1864
rect 22098 8900 22154 8936
rect 22098 8880 22100 8900
rect 22100 8880 22152 8900
rect 22152 8880 22154 8900
rect 22098 7384 22154 7440
rect 22098 6316 22154 6352
rect 22098 6296 22100 6316
rect 22100 6296 22152 6316
rect 22152 6296 22154 6316
rect 23294 30096 23350 30152
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 23386 29280 23442 29336
rect 23202 29028 23258 29064
rect 23202 29008 23204 29028
rect 23204 29008 23256 29028
rect 23256 29008 23258 29028
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 23386 27648 23442 27704
rect 22834 27376 22890 27432
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 23386 25916 23388 25936
rect 23388 25916 23440 25936
rect 23440 25916 23442 25936
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22742 21664 22798 21720
rect 23386 25880 23442 25916
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23202 20712 23258 20768
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22466 17060 22522 17096
rect 22466 17040 22468 17060
rect 22468 17040 22520 17060
rect 22520 17040 22522 17060
rect 22098 3052 22154 3088
rect 22098 3032 22100 3052
rect 22100 3032 22152 3052
rect 22152 3032 22154 3052
rect 23386 19488 23442 19544
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23386 18128 23442 18184
rect 24858 40704 24914 40760
rect 24306 36624 24362 36680
rect 24030 28464 24086 28520
rect 24674 38256 24730 38312
rect 24858 39888 24914 39944
rect 25318 39072 25374 39128
rect 24766 37440 24822 37496
rect 24490 34176 24546 34232
rect 24122 27276 24124 27296
rect 24124 27276 24176 27296
rect 24176 27276 24178 27296
rect 24122 27240 24178 27276
rect 23754 20576 23810 20632
rect 23662 20440 23718 20496
rect 25042 35808 25098 35864
rect 24582 27940 24638 27976
rect 24582 27920 24584 27940
rect 24584 27920 24636 27940
rect 24636 27920 24638 27940
rect 24950 27276 24952 27296
rect 24952 27276 25004 27296
rect 25004 27276 25006 27296
rect 24950 27240 25006 27276
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22926 17332 22982 17368
rect 22926 17312 22928 17332
rect 22928 17312 22980 17332
rect 22980 17312 22982 17332
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 23386 14592 23442 14648
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23294 12860 23296 12880
rect 23296 12860 23348 12880
rect 23348 12860 23350 12880
rect 23294 12824 23350 12860
rect 22282 3168 22338 3224
rect 22190 2352 22246 2408
rect 22282 1536 22338 1592
rect 22742 10512 22798 10568
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 23754 19624 23810 19680
rect 24030 19760 24086 19816
rect 23938 19372 23994 19408
rect 23938 19352 23940 19372
rect 23940 19352 23992 19372
rect 23992 19352 23994 19372
rect 23294 11600 23350 11656
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23202 10004 23204 10024
rect 23204 10004 23256 10024
rect 23256 10004 23258 10024
rect 23202 9968 23258 10004
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22650 4564 22652 4584
rect 22652 4564 22704 4584
rect 22704 4564 22706 4584
rect 22650 4528 22706 4564
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23386 4800 23442 4856
rect 23386 3984 23442 4040
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23938 13776 23994 13832
rect 24306 18808 24362 18864
rect 23938 12824 23994 12880
rect 23754 11756 23810 11792
rect 23754 11736 23756 11756
rect 23756 11736 23808 11756
rect 23808 11736 23810 11756
rect 23662 11192 23718 11248
rect 23294 1128 23350 1184
rect 23846 9868 23848 9888
rect 23848 9868 23900 9888
rect 23900 9868 23902 9888
rect 23846 9832 23902 9868
rect 23846 7268 23902 7304
rect 23846 7248 23848 7268
rect 23848 7248 23900 7268
rect 23900 7248 23902 7268
rect 24950 25220 25006 25256
rect 24950 25200 24952 25220
rect 24952 25200 25004 25220
rect 25004 25200 25006 25220
rect 24766 24384 24822 24440
rect 24490 23568 24546 23624
rect 24582 21936 24638 21992
rect 24858 23976 24914 24032
rect 24766 18672 24822 18728
rect 24582 17584 24638 17640
rect 24950 23704 25006 23760
rect 24950 22752 25006 22808
rect 25042 21936 25098 21992
rect 24950 21836 24952 21856
rect 24952 21836 25004 21856
rect 25004 21836 25006 21856
rect 24950 21800 25006 21836
rect 25410 22480 25466 22536
rect 24950 20304 25006 20360
rect 24858 17856 24914 17912
rect 24674 15136 24730 15192
rect 24582 13268 24584 13288
rect 24584 13268 24636 13288
rect 24636 13268 24638 13288
rect 24582 13232 24638 13268
rect 23938 5228 23994 5264
rect 23938 5208 23940 5228
rect 23940 5208 23992 5228
rect 23992 5208 23994 5228
rect 23846 3576 23902 3632
rect 24214 3732 24270 3768
rect 24214 3712 24216 3732
rect 24216 3712 24268 3732
rect 24268 3712 24270 3732
rect 24766 12960 24822 13016
rect 24858 12144 24914 12200
rect 24858 11328 24914 11384
rect 24766 10512 24822 10568
rect 24858 8880 24914 8936
rect 24858 8064 24914 8120
rect 24766 7248 24822 7304
rect 24674 6840 24730 6896
rect 24582 5616 24638 5672
rect 24766 5616 24822 5672
rect 25134 19252 25136 19272
rect 25136 19252 25188 19272
rect 25188 19252 25190 19272
rect 25134 19216 25190 19252
rect 25134 17040 25190 17096
rect 25042 16224 25098 16280
rect 25042 15428 25098 15464
rect 25042 15408 25044 15428
rect 25044 15408 25096 15428
rect 25096 15408 25098 15428
rect 25134 9696 25190 9752
rect 25042 6432 25098 6488
rect 25870 15272 25926 15328
rect 24950 720 25006 776
<< metal3 >>
rect 24117 56266 24183 56269
rect 26200 56266 27000 56296
rect 24117 56264 27000 56266
rect 24117 56208 24122 56264
rect 24178 56208 27000 56264
rect 24117 56206 27000 56208
rect 24117 56203 24183 56206
rect 26200 56176 27000 56206
rect 22369 55450 22435 55453
rect 26200 55450 27000 55480
rect 22369 55448 27000 55450
rect 22369 55392 22374 55448
rect 22430 55392 27000 55448
rect 22369 55390 27000 55392
rect 22369 55387 22435 55390
rect 26200 55360 27000 55390
rect 22829 54634 22895 54637
rect 26200 54634 27000 54664
rect 22829 54632 27000 54634
rect 22829 54576 22834 54632
rect 22890 54576 27000 54632
rect 22829 54574 27000 54576
rect 22829 54571 22895 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 23381 53818 23447 53821
rect 26200 53818 27000 53848
rect 23381 53816 27000 53818
rect 23381 53760 23386 53816
rect 23442 53760 27000 53816
rect 23381 53758 27000 53760
rect 23381 53755 23447 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 24577 53002 24643 53005
rect 26200 53002 27000 53032
rect 24577 53000 27000 53002
rect 24577 52944 24582 53000
rect 24638 52944 27000 53000
rect 24577 52942 27000 52944
rect 24577 52939 24643 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24945 52186 25011 52189
rect 26200 52186 27000 52216
rect 24945 52184 27000 52186
rect 24945 52128 24950 52184
rect 25006 52128 27000 52184
rect 24945 52126 27000 52128
rect 24945 52123 25011 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 24945 51370 25011 51373
rect 26200 51370 27000 51400
rect 24945 51368 27000 51370
rect 24945 51312 24950 51368
rect 25006 51312 27000 51368
rect 24945 51310 27000 51312
rect 24945 51307 25011 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 24945 50554 25011 50557
rect 26200 50554 27000 50584
rect 24945 50552 27000 50554
rect 24945 50496 24950 50552
rect 25006 50496 27000 50552
rect 24945 50494 27000 50496
rect 24945 50491 25011 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25497 49738 25563 49741
rect 26200 49738 27000 49768
rect 25497 49736 27000 49738
rect 25497 49680 25502 49736
rect 25558 49680 27000 49736
rect 25497 49678 27000 49680
rect 25497 49675 25563 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25129 48922 25195 48925
rect 26200 48922 27000 48952
rect 25129 48920 27000 48922
rect 25129 48864 25134 48920
rect 25190 48864 27000 48920
rect 25129 48862 27000 48864
rect 25129 48859 25195 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 25129 48106 25195 48109
rect 26200 48106 27000 48136
rect 25129 48104 27000 48106
rect 25129 48048 25134 48104
rect 25190 48048 27000 48104
rect 25129 48046 27000 48048
rect 25129 48043 25195 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 21030 47636 21036 47700
rect 21100 47698 21106 47700
rect 24761 47698 24827 47701
rect 21100 47696 24827 47698
rect 21100 47640 24766 47696
rect 24822 47640 24827 47696
rect 21100 47638 24827 47640
rect 21100 47636 21106 47638
rect 24761 47635 24827 47638
rect 16246 47500 16252 47564
rect 16316 47562 16322 47564
rect 25221 47562 25287 47565
rect 16316 47560 25287 47562
rect 16316 47504 25226 47560
rect 25282 47504 25287 47560
rect 16316 47502 25287 47504
rect 16316 47500 16322 47502
rect 25221 47499 25287 47502
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 20478 46956 20484 47020
rect 20548 47018 20554 47020
rect 24853 47018 24919 47021
rect 20548 47016 24919 47018
rect 20548 46960 24858 47016
rect 24914 46960 24919 47016
rect 20548 46958 24919 46960
rect 20548 46956 20554 46958
rect 24853 46955 24919 46958
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24761 44026 24827 44029
rect 26200 44026 27000 44056
rect 24761 44024 27000 44026
rect 24761 43968 24766 44024
rect 24822 43968 27000 44024
rect 24761 43966 27000 43968
rect 24761 43963 24827 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 25497 43210 25563 43213
rect 26200 43210 27000 43240
rect 25497 43208 27000 43210
rect 25497 43152 25502 43208
rect 25558 43152 27000 43208
rect 25497 43150 27000 43152
rect 25497 43147 25563 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 15326 42604 15332 42668
rect 15396 42666 15402 42668
rect 25221 42666 25287 42669
rect 15396 42664 25287 42666
rect 15396 42608 25226 42664
rect 25282 42608 25287 42664
rect 15396 42606 25287 42608
rect 15396 42604 15402 42606
rect 25221 42603 25287 42606
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25129 42394 25195 42397
rect 26200 42394 27000 42424
rect 25129 42392 27000 42394
rect 25129 42336 25134 42392
rect 25190 42336 27000 42392
rect 25129 42334 27000 42336
rect 25129 42331 25195 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 12198 41516 12204 41580
rect 12268 41578 12274 41580
rect 24853 41578 24919 41581
rect 12268 41576 24919 41578
rect 12268 41520 24858 41576
rect 24914 41520 24919 41576
rect 12268 41518 24919 41520
rect 12268 41516 12274 41518
rect 24853 41515 24919 41518
rect 25129 41578 25195 41581
rect 26200 41578 27000 41608
rect 25129 41576 27000 41578
rect 25129 41520 25134 41576
rect 25190 41520 27000 41576
rect 25129 41518 27000 41520
rect 25129 41515 25195 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 24853 40762 24919 40765
rect 26200 40762 27000 40792
rect 24853 40760 27000 40762
rect 24853 40704 24858 40760
rect 24914 40704 27000 40760
rect 24853 40702 27000 40704
rect 24853 40699 24919 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 19742 40020 19748 40084
rect 19812 40082 19818 40084
rect 23473 40082 23539 40085
rect 19812 40080 23539 40082
rect 19812 40024 23478 40080
rect 23534 40024 23539 40080
rect 19812 40022 23539 40024
rect 19812 40020 19818 40022
rect 23473 40019 23539 40022
rect 24853 39946 24919 39949
rect 26200 39946 27000 39976
rect 24853 39944 27000 39946
rect 24853 39888 24858 39944
rect 24914 39888 27000 39944
rect 24853 39886 27000 39888
rect 24853 39883 24919 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 24669 38314 24735 38317
rect 26200 38314 27000 38344
rect 24669 38312 27000 38314
rect 24669 38256 24674 38312
rect 24730 38256 27000 38312
rect 24669 38254 27000 38256
rect 24669 38251 24735 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 24761 37498 24827 37501
rect 26200 37498 27000 37528
rect 24761 37496 27000 37498
rect 24761 37440 24766 37496
rect 24822 37440 27000 37496
rect 24761 37438 27000 37440
rect 24761 37435 24827 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 24301 36682 24367 36685
rect 26200 36682 27000 36712
rect 24301 36680 27000 36682
rect 24301 36624 24306 36680
rect 24362 36624 27000 36680
rect 24301 36622 27000 36624
rect 24301 36619 24367 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 16430 35804 16436 35868
rect 16500 35866 16506 35868
rect 17033 35866 17099 35869
rect 16500 35864 17099 35866
rect 16500 35808 17038 35864
rect 17094 35808 17099 35864
rect 16500 35806 17099 35808
rect 16500 35804 16506 35806
rect 17033 35803 17099 35806
rect 25037 35866 25103 35869
rect 26200 35866 27000 35896
rect 25037 35864 27000 35866
rect 25037 35808 25042 35864
rect 25098 35808 27000 35864
rect 25037 35806 27000 35808
rect 25037 35803 25103 35806
rect 26200 35776 27000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 22737 35050 22803 35053
rect 26200 35050 27000 35080
rect 22737 35048 27000 35050
rect 22737 34992 22742 35048
rect 22798 34992 27000 35048
rect 22737 34990 27000 34992
rect 22737 34987 22803 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 15694 34444 15700 34508
rect 15764 34506 15770 34508
rect 17309 34506 17375 34509
rect 15764 34504 17375 34506
rect 15764 34448 17314 34504
rect 17370 34448 17375 34504
rect 15764 34446 17375 34448
rect 15764 34444 15770 34446
rect 17309 34443 17375 34446
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 24485 34234 24551 34237
rect 26200 34234 27000 34264
rect 24485 34232 27000 34234
rect 24485 34176 24490 34232
rect 24546 34176 27000 34232
rect 24485 34174 27000 34176
rect 24485 34171 24551 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 22093 33418 22159 33421
rect 26200 33418 27000 33448
rect 22093 33416 27000 33418
rect 22093 33360 22098 33416
rect 22154 33360 27000 33416
rect 22093 33358 27000 33360
rect 22093 33355 22159 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 21817 32602 21883 32605
rect 26200 32602 27000 32632
rect 21817 32600 27000 32602
rect 21817 32544 21822 32600
rect 21878 32544 27000 32600
rect 21817 32542 27000 32544
rect 21817 32539 21883 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 22093 31786 22159 31789
rect 26200 31786 27000 31816
rect 22093 31784 27000 31786
rect 22093 31728 22098 31784
rect 22154 31728 27000 31784
rect 22093 31726 27000 31728
rect 22093 31723 22159 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 22093 31242 22159 31245
rect 22093 31240 23490 31242
rect 22093 31184 22098 31240
rect 22154 31184 23490 31240
rect 22093 31182 23490 31184
rect 22093 31179 22159 31182
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 23430 30970 23490 31182
rect 26200 30970 27000 31000
rect 23430 30910 27000 30970
rect 26200 30880 27000 30910
rect 18597 30836 18663 30837
rect 18597 30834 18644 30836
rect 18552 30832 18644 30834
rect 18552 30776 18602 30832
rect 18552 30774 18644 30776
rect 18597 30772 18644 30774
rect 18708 30772 18714 30836
rect 18597 30771 18663 30772
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 23289 30154 23355 30157
rect 26200 30154 27000 30184
rect 23289 30152 27000 30154
rect 23289 30096 23294 30152
rect 23350 30096 27000 30152
rect 23289 30094 27000 30096
rect 23289 30091 23355 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 12709 29746 12775 29749
rect 15285 29746 15351 29749
rect 12709 29744 15351 29746
rect 12709 29688 12714 29744
rect 12770 29688 15290 29744
rect 15346 29688 15351 29744
rect 12709 29686 15351 29688
rect 12709 29683 12775 29686
rect 15285 29683 15351 29686
rect 13537 29610 13603 29613
rect 18689 29610 18755 29613
rect 13537 29608 18755 29610
rect 13537 29552 13542 29608
rect 13598 29552 18694 29608
rect 18750 29552 18755 29608
rect 13537 29550 18755 29552
rect 13537 29547 13603 29550
rect 18689 29547 18755 29550
rect 10133 29474 10199 29477
rect 12985 29474 13051 29477
rect 16021 29474 16087 29477
rect 10133 29472 16087 29474
rect 10133 29416 10138 29472
rect 10194 29416 12990 29472
rect 13046 29416 16026 29472
rect 16082 29416 16087 29472
rect 10133 29414 16087 29416
rect 10133 29411 10199 29414
rect 12985 29411 13051 29414
rect 16021 29411 16087 29414
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 13813 29338 13879 29341
rect 15101 29338 15167 29341
rect 13813 29336 15167 29338
rect 13813 29280 13818 29336
rect 13874 29280 15106 29336
rect 15162 29280 15167 29336
rect 13813 29278 15167 29280
rect 13813 29275 13879 29278
rect 15101 29275 15167 29278
rect 23381 29338 23447 29341
rect 26200 29338 27000 29368
rect 23381 29336 27000 29338
rect 23381 29280 23386 29336
rect 23442 29280 27000 29336
rect 23381 29278 27000 29280
rect 23381 29275 23447 29278
rect 26200 29248 27000 29278
rect 13721 29202 13787 29205
rect 19057 29202 19123 29205
rect 13721 29200 19123 29202
rect 13721 29144 13726 29200
rect 13782 29144 19062 29200
rect 19118 29144 19123 29200
rect 13721 29142 19123 29144
rect 13721 29139 13787 29142
rect 19057 29139 19123 29142
rect 4337 29066 4403 29069
rect 22001 29066 22067 29069
rect 4337 29064 22067 29066
rect 4337 29008 4342 29064
rect 4398 29008 22006 29064
rect 22062 29008 22067 29064
rect 4337 29006 22067 29008
rect 4337 29003 4403 29006
rect 22001 29003 22067 29006
rect 22686 29004 22692 29068
rect 22756 29066 22762 29068
rect 23197 29066 23263 29069
rect 22756 29064 23263 29066
rect 22756 29008 23202 29064
rect 23258 29008 23263 29064
rect 22756 29006 23263 29008
rect 22756 29004 22762 29006
rect 23197 29003 23263 29006
rect 15653 28930 15719 28933
rect 17493 28930 17559 28933
rect 15653 28928 17559 28930
rect 15653 28872 15658 28928
rect 15714 28872 17498 28928
rect 17554 28872 17559 28928
rect 15653 28870 17559 28872
rect 15653 28867 15719 28870
rect 17493 28867 17559 28870
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 15285 28658 15351 28661
rect 15929 28658 15995 28661
rect 15285 28656 15995 28658
rect 15285 28600 15290 28656
rect 15346 28600 15934 28656
rect 15990 28600 15995 28656
rect 15285 28598 15995 28600
rect 15285 28595 15351 28598
rect 15929 28595 15995 28598
rect 24025 28522 24091 28525
rect 26200 28522 27000 28552
rect 24025 28520 27000 28522
rect 24025 28464 24030 28520
rect 24086 28464 27000 28520
rect 24025 28462 27000 28464
rect 24025 28459 24091 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 10961 27978 11027 27981
rect 24577 27978 24643 27981
rect 10961 27976 24643 27978
rect 10961 27920 10966 27976
rect 11022 27920 24582 27976
rect 24638 27920 24643 27976
rect 10961 27918 24643 27920
rect 10961 27915 11027 27918
rect 24577 27915 24643 27918
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 23381 27706 23447 27709
rect 26200 27706 27000 27736
rect 23381 27704 27000 27706
rect 23381 27648 23386 27704
rect 23442 27648 27000 27704
rect 23381 27646 27000 27648
rect 23381 27643 23447 27646
rect 26200 27616 27000 27646
rect 18638 27508 18644 27572
rect 18708 27570 18714 27572
rect 18781 27570 18847 27573
rect 18708 27568 18847 27570
rect 18708 27512 18786 27568
rect 18842 27512 18847 27568
rect 18708 27510 18847 27512
rect 18708 27508 18714 27510
rect 18781 27507 18847 27510
rect 5533 27434 5599 27437
rect 22829 27434 22895 27437
rect 5533 27432 22895 27434
rect 5533 27376 5538 27432
rect 5594 27376 22834 27432
rect 22890 27376 22895 27432
rect 5533 27374 22895 27376
rect 5533 27371 5599 27374
rect 22829 27371 22895 27374
rect 9305 27298 9371 27301
rect 14457 27298 14523 27301
rect 9305 27296 14523 27298
rect 9305 27240 9310 27296
rect 9366 27240 14462 27296
rect 14518 27240 14523 27296
rect 9305 27238 14523 27240
rect 9305 27235 9371 27238
rect 14457 27235 14523 27238
rect 14733 27298 14799 27301
rect 16297 27298 16363 27301
rect 14733 27296 16363 27298
rect 14733 27240 14738 27296
rect 14794 27240 16302 27296
rect 16358 27240 16363 27296
rect 14733 27238 16363 27240
rect 14733 27235 14799 27238
rect 16297 27235 16363 27238
rect 24117 27298 24183 27301
rect 24945 27298 25011 27301
rect 24117 27296 25011 27298
rect 24117 27240 24122 27296
rect 24178 27240 24950 27296
rect 25006 27240 25011 27296
rect 24117 27238 25011 27240
rect 24117 27235 24183 27238
rect 24945 27235 25011 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 22277 26890 22343 26893
rect 26200 26890 27000 26920
rect 22277 26888 27000 26890
rect 22277 26832 22282 26888
rect 22338 26832 27000 26888
rect 22277 26830 27000 26832
rect 22277 26827 22343 26830
rect 26200 26800 27000 26830
rect 13721 26754 13787 26757
rect 22461 26754 22527 26757
rect 13721 26752 22527 26754
rect 13721 26696 13726 26752
rect 13782 26696 22466 26752
rect 22522 26696 22527 26752
rect 13721 26694 22527 26696
rect 13721 26691 13787 26694
rect 22461 26691 22527 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 10317 26482 10383 26485
rect 17125 26482 17191 26485
rect 10317 26480 17191 26482
rect 10317 26424 10322 26480
rect 10378 26424 17130 26480
rect 17186 26424 17191 26480
rect 10317 26422 17191 26424
rect 10317 26419 10383 26422
rect 17125 26419 17191 26422
rect 17718 26420 17724 26484
rect 17788 26482 17794 26484
rect 18689 26482 18755 26485
rect 17788 26480 18755 26482
rect 17788 26424 18694 26480
rect 18750 26424 18755 26480
rect 17788 26422 18755 26424
rect 17788 26420 17794 26422
rect 18689 26419 18755 26422
rect 18965 26348 19031 26349
rect 18965 26346 19012 26348
rect 18920 26344 19012 26346
rect 18920 26288 18970 26344
rect 18920 26286 19012 26288
rect 18965 26284 19012 26286
rect 19076 26284 19082 26348
rect 18965 26283 19031 26284
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 10593 26074 10659 26077
rect 22369 26074 22435 26077
rect 26200 26074 27000 26104
rect 10593 26072 12450 26074
rect 10593 26016 10598 26072
rect 10654 26016 12450 26072
rect 10593 26014 12450 26016
rect 10593 26011 10659 26014
rect 12390 25938 12450 26014
rect 22369 26072 27000 26074
rect 22369 26016 22374 26072
rect 22430 26016 27000 26072
rect 22369 26014 27000 26016
rect 22369 26011 22435 26014
rect 26200 25984 27000 26014
rect 23381 25938 23447 25941
rect 12390 25936 23447 25938
rect 12390 25880 23386 25936
rect 23442 25880 23447 25936
rect 12390 25878 23447 25880
rect 23381 25875 23447 25878
rect 11646 25740 11652 25804
rect 11716 25802 11722 25804
rect 18045 25802 18111 25805
rect 11716 25800 18111 25802
rect 11716 25744 18050 25800
rect 18106 25744 18111 25800
rect 11716 25742 18111 25744
rect 11716 25740 11722 25742
rect 18045 25739 18111 25742
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 14457 25530 14523 25533
rect 14457 25528 22110 25530
rect 14457 25472 14462 25528
rect 14518 25472 22110 25528
rect 14457 25470 22110 25472
rect 14457 25467 14523 25470
rect 16113 25394 16179 25397
rect 16246 25394 16252 25396
rect 16113 25392 16252 25394
rect 16113 25336 16118 25392
rect 16174 25336 16252 25392
rect 16113 25334 16252 25336
rect 16113 25331 16179 25334
rect 16246 25332 16252 25334
rect 16316 25332 16322 25396
rect 20713 25394 20779 25397
rect 21030 25394 21036 25396
rect 20713 25392 21036 25394
rect 20713 25336 20718 25392
rect 20774 25336 21036 25392
rect 20713 25334 21036 25336
rect 20713 25331 20779 25334
rect 21030 25332 21036 25334
rect 21100 25332 21106 25396
rect 22050 25394 22110 25470
rect 24710 25394 24716 25396
rect 22050 25334 24716 25394
rect 24710 25332 24716 25334
rect 24780 25332 24786 25396
rect 24945 25258 25011 25261
rect 26200 25258 27000 25288
rect 24945 25256 27000 25258
rect 24945 25200 24950 25256
rect 25006 25200 27000 25256
rect 24945 25198 27000 25200
rect 24945 25195 25011 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 20805 24988 20871 24989
rect 20805 24984 20852 24988
rect 20916 24986 20922 24988
rect 21817 24986 21883 24989
rect 22134 24986 22140 24988
rect 20805 24928 20810 24984
rect 20805 24924 20852 24928
rect 20916 24926 20962 24986
rect 21817 24984 22140 24986
rect 21817 24928 21822 24984
rect 21878 24928 22140 24984
rect 21817 24926 22140 24928
rect 20916 24924 20922 24926
rect 20805 24923 20871 24924
rect 21817 24923 21883 24926
rect 22134 24924 22140 24926
rect 22204 24924 22210 24988
rect 8937 24714 9003 24717
rect 18505 24714 18571 24717
rect 8937 24712 18571 24714
rect 8937 24656 8942 24712
rect 8998 24656 18510 24712
rect 18566 24656 18571 24712
rect 8937 24654 18571 24656
rect 8937 24651 9003 24654
rect 18505 24651 18571 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24761 24442 24827 24445
rect 26200 24442 27000 24472
rect 24761 24440 27000 24442
rect 24761 24384 24766 24440
rect 24822 24384 27000 24440
rect 24761 24382 27000 24384
rect 24761 24379 24827 24382
rect 26200 24352 27000 24382
rect 12617 24170 12683 24173
rect 14825 24170 14891 24173
rect 12617 24168 14891 24170
rect 12617 24112 12622 24168
rect 12678 24112 14830 24168
rect 14886 24112 14891 24168
rect 12617 24110 14891 24112
rect 12617 24107 12683 24110
rect 14825 24107 14891 24110
rect 13445 24034 13511 24037
rect 14641 24034 14707 24037
rect 13445 24032 14707 24034
rect 13445 23976 13450 24032
rect 13506 23976 14646 24032
rect 14702 23976 14707 24032
rect 13445 23974 14707 23976
rect 13445 23971 13511 23974
rect 14641 23971 14707 23974
rect 20437 24034 20503 24037
rect 24853 24034 24919 24037
rect 20437 24032 24919 24034
rect 20437 23976 20442 24032
rect 20498 23976 24858 24032
rect 24914 23976 24919 24032
rect 20437 23974 24919 23976
rect 20437 23971 20503 23974
rect 24853 23971 24919 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 13261 23898 13327 23901
rect 13261 23896 16682 23898
rect 13261 23840 13266 23896
rect 13322 23840 16682 23896
rect 13261 23838 16682 23840
rect 13261 23835 13327 23838
rect 13997 23762 14063 23765
rect 16481 23762 16547 23765
rect 13997 23760 16547 23762
rect 13997 23704 14002 23760
rect 14058 23704 16486 23760
rect 16542 23704 16547 23760
rect 13997 23702 16547 23704
rect 16622 23762 16682 23838
rect 24945 23762 25011 23765
rect 16622 23760 25011 23762
rect 16622 23704 24950 23760
rect 25006 23704 25011 23760
rect 16622 23702 25011 23704
rect 13997 23699 14063 23702
rect 16481 23699 16547 23702
rect 24945 23699 25011 23702
rect 7189 23626 7255 23629
rect 16389 23626 16455 23629
rect 22001 23626 22067 23629
rect 7189 23624 16455 23626
rect 7189 23568 7194 23624
rect 7250 23568 16394 23624
rect 16450 23568 16455 23624
rect 7189 23566 16455 23568
rect 7189 23563 7255 23566
rect 16389 23563 16455 23566
rect 16622 23624 22067 23626
rect 16622 23568 22006 23624
rect 22062 23568 22067 23624
rect 16622 23566 22067 23568
rect 13486 23428 13492 23492
rect 13556 23490 13562 23492
rect 14273 23490 14339 23493
rect 13556 23488 14339 23490
rect 13556 23432 14278 23488
rect 14334 23432 14339 23488
rect 13556 23430 14339 23432
rect 13556 23428 13562 23430
rect 14273 23427 14339 23430
rect 15101 23490 15167 23493
rect 16622 23490 16682 23566
rect 22001 23563 22067 23566
rect 24485 23626 24551 23629
rect 26200 23626 27000 23656
rect 24485 23624 27000 23626
rect 24485 23568 24490 23624
rect 24546 23568 27000 23624
rect 24485 23566 27000 23568
rect 24485 23563 24551 23566
rect 26200 23536 27000 23566
rect 15101 23488 16682 23490
rect 15101 23432 15106 23488
rect 15162 23432 16682 23488
rect 15101 23430 16682 23432
rect 19517 23490 19583 23493
rect 20989 23490 21055 23493
rect 19517 23488 21055 23490
rect 19517 23432 19522 23488
rect 19578 23432 20994 23488
rect 21050 23432 21055 23488
rect 19517 23430 21055 23432
rect 15101 23427 15167 23430
rect 19517 23427 19583 23430
rect 20989 23427 21055 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 6269 23218 6335 23221
rect 22093 23218 22159 23221
rect 6269 23216 22159 23218
rect 6269 23160 6274 23216
rect 6330 23160 22098 23216
rect 22154 23160 22159 23216
rect 6269 23158 22159 23160
rect 6269 23155 6335 23158
rect 22093 23155 22159 23158
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 24945 22810 25011 22813
rect 26200 22810 27000 22840
rect 24945 22808 27000 22810
rect 24945 22752 24950 22808
rect 25006 22752 27000 22808
rect 24945 22750 27000 22752
rect 24945 22747 25011 22750
rect 26200 22720 27000 22750
rect 16389 22674 16455 22677
rect 24526 22674 24532 22676
rect 16389 22672 24532 22674
rect 16389 22616 16394 22672
rect 16450 22616 24532 22672
rect 16389 22614 24532 22616
rect 16389 22611 16455 22614
rect 24526 22612 24532 22614
rect 24596 22612 24602 22676
rect 10910 22476 10916 22540
rect 10980 22538 10986 22540
rect 16389 22538 16455 22541
rect 10980 22536 16455 22538
rect 10980 22480 16394 22536
rect 16450 22480 16455 22536
rect 10980 22478 16455 22480
rect 10980 22476 10986 22478
rect 16389 22475 16455 22478
rect 18781 22538 18847 22541
rect 25405 22538 25471 22541
rect 18781 22536 25471 22538
rect 18781 22480 18786 22536
rect 18842 22480 25410 22536
rect 25466 22480 25471 22536
rect 18781 22478 25471 22480
rect 18781 22475 18847 22478
rect 25405 22475 25471 22478
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 9121 22130 9187 22133
rect 21909 22130 21975 22133
rect 9121 22128 21975 22130
rect 9121 22072 9126 22128
rect 9182 22072 21914 22128
rect 21970 22072 21975 22128
rect 9121 22070 21975 22072
rect 9121 22067 9187 22070
rect 21909 22067 21975 22070
rect 6545 21994 6611 21997
rect 24577 21994 24643 21997
rect 6545 21992 24643 21994
rect 6545 21936 6550 21992
rect 6606 21936 24582 21992
rect 24638 21936 24643 21992
rect 6545 21934 24643 21936
rect 6545 21931 6611 21934
rect 24577 21931 24643 21934
rect 25037 21994 25103 21997
rect 26200 21994 27000 22024
rect 25037 21992 27000 21994
rect 25037 21936 25042 21992
rect 25098 21936 27000 21992
rect 25037 21934 27000 21936
rect 25037 21931 25103 21934
rect 26200 21904 27000 21934
rect 19333 21858 19399 21861
rect 19609 21858 19675 21861
rect 19333 21856 19675 21858
rect 19333 21800 19338 21856
rect 19394 21800 19614 21856
rect 19670 21800 19675 21856
rect 19333 21798 19675 21800
rect 19333 21795 19399 21798
rect 19609 21795 19675 21798
rect 21909 21858 21975 21861
rect 24945 21858 25011 21861
rect 21909 21856 25011 21858
rect 21909 21800 21914 21856
rect 21970 21800 24950 21856
rect 25006 21800 25011 21856
rect 21909 21798 25011 21800
rect 21909 21795 21975 21798
rect 24945 21795 25011 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 22001 21722 22067 21725
rect 22737 21722 22803 21725
rect 22001 21720 22803 21722
rect 22001 21664 22006 21720
rect 22062 21664 22742 21720
rect 22798 21664 22803 21720
rect 22001 21662 22803 21664
rect 22001 21659 22067 21662
rect 22737 21659 22803 21662
rect 4654 21524 4660 21588
rect 4724 21586 4730 21588
rect 22185 21586 22251 21589
rect 4724 21584 22251 21586
rect 4724 21528 22190 21584
rect 22246 21528 22251 21584
rect 4724 21526 22251 21528
rect 4724 21524 4730 21526
rect 22185 21523 22251 21526
rect 5165 21450 5231 21453
rect 16389 21450 16455 21453
rect 5165 21448 16455 21450
rect 5165 21392 5170 21448
rect 5226 21392 16394 21448
rect 16450 21392 16455 21448
rect 5165 21390 16455 21392
rect 5165 21387 5231 21390
rect 16389 21387 16455 21390
rect 17125 21450 17191 21453
rect 20478 21450 20484 21452
rect 17125 21448 20484 21450
rect 17125 21392 17130 21448
rect 17186 21392 20484 21448
rect 17125 21390 20484 21392
rect 17125 21387 17191 21390
rect 20478 21388 20484 21390
rect 20548 21388 20554 21452
rect 22461 21450 22527 21453
rect 22461 21448 24042 21450
rect 22461 21392 22466 21448
rect 22522 21392 24042 21448
rect 22461 21390 24042 21392
rect 22461 21387 22527 21390
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 13629 21178 13695 21181
rect 17534 21178 17540 21180
rect 13629 21176 17540 21178
rect 13629 21120 13634 21176
rect 13690 21120 17540 21176
rect 13629 21118 17540 21120
rect 13629 21115 13695 21118
rect 17534 21116 17540 21118
rect 17604 21116 17610 21180
rect 23982 21178 24042 21390
rect 26200 21178 27000 21208
rect 23982 21118 27000 21178
rect 26200 21088 27000 21118
rect 19333 21042 19399 21045
rect 12390 21040 19399 21042
rect 12390 20984 19338 21040
rect 19394 20984 19399 21040
rect 12390 20982 19399 20984
rect 12390 20906 12450 20982
rect 19333 20979 19399 20982
rect 6686 20846 12450 20906
rect 6686 20501 6746 20846
rect 12566 20844 12572 20908
rect 12636 20906 12642 20908
rect 19425 20906 19491 20909
rect 12636 20904 19491 20906
rect 12636 20848 19430 20904
rect 19486 20848 19491 20904
rect 12636 20846 19491 20848
rect 12636 20844 12642 20846
rect 19425 20843 19491 20846
rect 21265 20906 21331 20909
rect 21817 20906 21883 20909
rect 21265 20904 21883 20906
rect 21265 20848 21270 20904
rect 21326 20848 21822 20904
rect 21878 20848 21883 20904
rect 21265 20846 21883 20848
rect 21265 20843 21331 20846
rect 21817 20843 21883 20846
rect 14181 20772 14247 20773
rect 14181 20768 14228 20772
rect 14292 20770 14298 20772
rect 20805 20770 20871 20773
rect 23197 20770 23263 20773
rect 14181 20712 14186 20768
rect 14181 20708 14228 20712
rect 14292 20710 14338 20770
rect 20805 20768 23263 20770
rect 20805 20712 20810 20768
rect 20866 20712 23202 20768
rect 23258 20712 23263 20768
rect 20805 20710 23263 20712
rect 14292 20708 14298 20710
rect 14181 20707 14247 20708
rect 20805 20707 20871 20710
rect 23197 20707 23263 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 11973 20634 12039 20637
rect 14825 20634 14891 20637
rect 11973 20632 14891 20634
rect 11973 20576 11978 20632
rect 12034 20576 14830 20632
rect 14886 20576 14891 20632
rect 11973 20574 14891 20576
rect 11973 20571 12039 20574
rect 14825 20571 14891 20574
rect 17493 20634 17559 20637
rect 17677 20634 17743 20637
rect 23749 20634 23815 20637
rect 17493 20632 17743 20634
rect 17493 20576 17498 20632
rect 17554 20576 17682 20632
rect 17738 20576 17743 20632
rect 17493 20574 17743 20576
rect 17493 20571 17559 20574
rect 17677 20571 17743 20574
rect 18462 20632 23815 20634
rect 18462 20576 23754 20632
rect 23810 20576 23815 20632
rect 18462 20574 23815 20576
rect 6686 20496 6795 20501
rect 6686 20440 6734 20496
rect 6790 20440 6795 20496
rect 6686 20438 6795 20440
rect 6729 20435 6795 20438
rect 8109 20498 8175 20501
rect 18462 20498 18522 20574
rect 23749 20571 23815 20574
rect 8109 20496 18522 20498
rect 8109 20440 8114 20496
rect 8170 20440 18522 20496
rect 8109 20438 18522 20440
rect 18965 20498 19031 20501
rect 23657 20498 23723 20501
rect 18965 20496 23723 20498
rect 18965 20440 18970 20496
rect 19026 20440 23662 20496
rect 23718 20440 23723 20496
rect 18965 20438 23723 20440
rect 8109 20435 8175 20438
rect 18965 20435 19031 20438
rect 23657 20435 23723 20438
rect 8385 20362 8451 20365
rect 22001 20362 22067 20365
rect 8385 20360 22067 20362
rect 8385 20304 8390 20360
rect 8446 20304 22006 20360
rect 22062 20304 22067 20360
rect 8385 20302 22067 20304
rect 8385 20299 8451 20302
rect 22001 20299 22067 20302
rect 24945 20362 25011 20365
rect 26200 20362 27000 20392
rect 24945 20360 27000 20362
rect 24945 20304 24950 20360
rect 25006 20304 27000 20360
rect 24945 20302 27000 20304
rect 24945 20299 25011 20302
rect 26200 20272 27000 20302
rect 7373 20226 7439 20229
rect 12433 20226 12499 20229
rect 7373 20224 12499 20226
rect 7373 20168 7378 20224
rect 7434 20168 12438 20224
rect 12494 20168 12499 20224
rect 7373 20166 12499 20168
rect 7373 20163 7439 20166
rect 12433 20163 12499 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 5349 20090 5415 20093
rect 8661 20090 8727 20093
rect 5349 20088 8727 20090
rect 5349 20032 5354 20088
rect 5410 20032 8666 20088
rect 8722 20032 8727 20088
rect 5349 20030 8727 20032
rect 5349 20027 5415 20030
rect 8661 20027 8727 20030
rect 14365 20090 14431 20093
rect 18321 20090 18387 20093
rect 14365 20088 18387 20090
rect 14365 20032 14370 20088
rect 14426 20032 18326 20088
rect 18382 20032 18387 20088
rect 14365 20030 18387 20032
rect 14365 20027 14431 20030
rect 18321 20027 18387 20030
rect 3969 19954 4035 19957
rect 20805 19954 20871 19957
rect 3969 19952 20871 19954
rect 3969 19896 3974 19952
rect 4030 19896 20810 19952
rect 20866 19896 20871 19952
rect 3969 19894 20871 19896
rect 3969 19891 4035 19894
rect 20805 19891 20871 19894
rect 4613 19818 4679 19821
rect 8661 19818 8727 19821
rect 17585 19818 17651 19821
rect 4613 19816 8586 19818
rect 4613 19760 4618 19816
rect 4674 19760 8586 19816
rect 4613 19758 8586 19760
rect 4613 19755 4679 19758
rect 8526 19682 8586 19758
rect 8661 19816 17651 19818
rect 8661 19760 8666 19816
rect 8722 19760 17590 19816
rect 17646 19760 17651 19816
rect 8661 19758 17651 19760
rect 8661 19755 8727 19758
rect 17585 19755 17651 19758
rect 20713 19818 20779 19821
rect 24025 19818 24091 19821
rect 20713 19816 24091 19818
rect 20713 19760 20718 19816
rect 20774 19760 24030 19816
rect 24086 19760 24091 19816
rect 20713 19758 24091 19760
rect 20713 19755 20779 19758
rect 24025 19755 24091 19758
rect 20621 19684 20687 19685
rect 14958 19682 14964 19684
rect 8526 19622 14964 19682
rect 14958 19620 14964 19622
rect 15028 19620 15034 19684
rect 20621 19682 20668 19684
rect 20540 19680 20668 19682
rect 20732 19682 20738 19684
rect 23749 19682 23815 19685
rect 20732 19680 23815 19682
rect 20540 19624 20626 19680
rect 20732 19624 23754 19680
rect 23810 19624 23815 19680
rect 20540 19622 20668 19624
rect 20621 19620 20668 19622
rect 20732 19622 23815 19624
rect 20732 19620 20738 19622
rect 20621 19619 20687 19620
rect 23749 19619 23815 19622
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 9029 19546 9095 19549
rect 14549 19546 14615 19549
rect 9029 19544 14615 19546
rect 9029 19488 9034 19544
rect 9090 19488 14554 19544
rect 14610 19488 14615 19544
rect 9029 19486 14615 19488
rect 9029 19483 9095 19486
rect 14549 19483 14615 19486
rect 23381 19546 23447 19549
rect 26200 19546 27000 19576
rect 23381 19544 27000 19546
rect 23381 19488 23386 19544
rect 23442 19488 27000 19544
rect 23381 19486 27000 19488
rect 23381 19483 23447 19486
rect 26200 19456 27000 19486
rect 5073 19410 5139 19413
rect 15142 19410 15148 19412
rect 5073 19408 15148 19410
rect 5073 19352 5078 19408
rect 5134 19352 15148 19408
rect 5073 19350 15148 19352
rect 5073 19347 5139 19350
rect 15142 19348 15148 19350
rect 15212 19348 15218 19412
rect 17033 19410 17099 19413
rect 23933 19410 23999 19413
rect 17033 19408 23999 19410
rect 17033 19352 17038 19408
rect 17094 19352 23938 19408
rect 23994 19352 23999 19408
rect 17033 19350 23999 19352
rect 17033 19347 17099 19350
rect 23933 19347 23999 19350
rect 6177 19274 6243 19277
rect 25129 19274 25195 19277
rect 6177 19272 25195 19274
rect 6177 19216 6182 19272
rect 6238 19216 25134 19272
rect 25190 19216 25195 19272
rect 6177 19214 25195 19216
rect 6177 19211 6243 19214
rect 25129 19211 25195 19214
rect 15285 19138 15351 19141
rect 16982 19138 16988 19140
rect 15285 19136 16988 19138
rect 15285 19080 15290 19136
rect 15346 19080 16988 19136
rect 15285 19078 16988 19080
rect 15285 19075 15351 19078
rect 16982 19076 16988 19078
rect 17052 19076 17058 19140
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 14958 18940 14964 19004
rect 15028 19002 15034 19004
rect 21030 19002 21036 19004
rect 15028 18942 21036 19002
rect 15028 18940 15034 18942
rect 21030 18940 21036 18942
rect 21100 18940 21106 19004
rect 5717 18866 5783 18869
rect 5717 18864 12450 18866
rect 5717 18808 5722 18864
rect 5778 18808 12450 18864
rect 5717 18806 12450 18808
rect 5717 18803 5783 18806
rect 4061 18730 4127 18733
rect 12390 18730 12450 18806
rect 15142 18804 15148 18868
rect 15212 18866 15218 18868
rect 24301 18866 24367 18869
rect 15212 18864 24367 18866
rect 15212 18808 24306 18864
rect 24362 18808 24367 18864
rect 15212 18806 24367 18808
rect 15212 18804 15218 18806
rect 24301 18803 24367 18806
rect 20805 18730 20871 18733
rect 4061 18728 8402 18730
rect 4061 18672 4066 18728
rect 4122 18672 8402 18728
rect 4061 18670 8402 18672
rect 12390 18728 20871 18730
rect 12390 18672 20810 18728
rect 20866 18672 20871 18728
rect 12390 18670 20871 18672
rect 4061 18667 4127 18670
rect 8342 18594 8402 18670
rect 20805 18667 20871 18670
rect 24761 18730 24827 18733
rect 26200 18730 27000 18760
rect 24761 18728 27000 18730
rect 24761 18672 24766 18728
rect 24822 18672 27000 18728
rect 24761 18670 27000 18672
rect 24761 18667 24827 18670
rect 26200 18640 27000 18670
rect 15101 18594 15167 18597
rect 8342 18592 15167 18594
rect 8342 18536 15106 18592
rect 15162 18536 15167 18592
rect 8342 18534 15167 18536
rect 15101 18531 15167 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 9949 18458 10015 18461
rect 9446 18456 10015 18458
rect 9446 18400 9954 18456
rect 10010 18400 10015 18456
rect 9446 18398 10015 18400
rect 3550 18260 3556 18324
rect 3620 18322 3626 18324
rect 9446 18322 9506 18398
rect 9949 18395 10015 18398
rect 3620 18262 9506 18322
rect 9673 18322 9739 18325
rect 21909 18322 21975 18325
rect 9673 18320 21975 18322
rect 9673 18264 9678 18320
rect 9734 18264 21914 18320
rect 21970 18264 21975 18320
rect 9673 18262 21975 18264
rect 3620 18260 3626 18262
rect 9673 18259 9739 18262
rect 21909 18259 21975 18262
rect 4705 18186 4771 18189
rect 23381 18186 23447 18189
rect 4705 18184 23447 18186
rect 4705 18128 4710 18184
rect 4766 18128 23386 18184
rect 23442 18128 23447 18184
rect 4705 18126 23447 18128
rect 4705 18123 4771 18126
rect 23381 18123 23447 18126
rect 9213 18052 9279 18053
rect 11789 18052 11855 18053
rect 11973 18052 12039 18053
rect 9213 18048 9260 18052
rect 9324 18050 9330 18052
rect 11789 18050 11836 18052
rect 9213 17992 9218 18048
rect 9213 17988 9260 17992
rect 9324 17990 9370 18050
rect 11744 18048 11836 18050
rect 11744 17992 11794 18048
rect 11744 17990 11836 17992
rect 9324 17988 9330 17990
rect 11789 17988 11836 17990
rect 11900 17988 11906 18052
rect 11973 18048 12020 18052
rect 12084 18050 12090 18052
rect 11973 17992 11978 18048
rect 11973 17988 12020 17992
rect 12084 17990 12130 18050
rect 12084 17988 12090 17990
rect 14038 17988 14044 18052
rect 14108 18050 14114 18052
rect 14181 18050 14247 18053
rect 14108 18048 14247 18050
rect 14108 17992 14186 18048
rect 14242 17992 14247 18048
rect 14108 17990 14247 17992
rect 14108 17988 14114 17990
rect 9213 17987 9279 17988
rect 11789 17987 11855 17988
rect 11973 17987 12039 17988
rect 14181 17987 14247 17990
rect 15878 17988 15884 18052
rect 15948 18050 15954 18052
rect 16297 18050 16363 18053
rect 15948 18048 16363 18050
rect 15948 17992 16302 18048
rect 16358 17992 16363 18048
rect 15948 17990 16363 17992
rect 15948 17988 15954 17990
rect 16297 17987 16363 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 4521 17914 4587 17917
rect 15745 17916 15811 17917
rect 4521 17912 10058 17914
rect 4521 17856 4526 17912
rect 4582 17856 10058 17912
rect 4521 17854 10058 17856
rect 4521 17851 4587 17854
rect 1301 17778 1367 17781
rect 9765 17778 9831 17781
rect 1301 17776 9831 17778
rect 1301 17720 1306 17776
rect 1362 17720 9770 17776
rect 9826 17720 9831 17776
rect 1301 17718 9831 17720
rect 1301 17715 1367 17718
rect 9765 17715 9831 17718
rect 6085 17642 6151 17645
rect 9998 17642 10058 17854
rect 15694 17852 15700 17916
rect 15764 17914 15811 17916
rect 18781 17914 18847 17917
rect 22318 17914 22324 17916
rect 15764 17912 15856 17914
rect 15806 17856 15856 17912
rect 15764 17854 15856 17856
rect 18781 17912 22324 17914
rect 18781 17856 18786 17912
rect 18842 17856 22324 17912
rect 18781 17854 22324 17856
rect 15764 17852 15811 17854
rect 15745 17851 15811 17852
rect 18781 17851 18847 17854
rect 22318 17852 22324 17854
rect 22388 17852 22394 17916
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 10133 17778 10199 17781
rect 19057 17778 19123 17781
rect 10133 17776 19123 17778
rect 10133 17720 10138 17776
rect 10194 17720 19062 17776
rect 19118 17720 19123 17776
rect 10133 17718 19123 17720
rect 10133 17715 10199 17718
rect 19057 17715 19123 17718
rect 24577 17642 24643 17645
rect 6085 17640 8402 17642
rect 6085 17584 6090 17640
rect 6146 17584 8402 17640
rect 6085 17582 8402 17584
rect 9998 17640 24643 17642
rect 9998 17584 24582 17640
rect 24638 17584 24643 17640
rect 9998 17582 24643 17584
rect 6085 17579 6151 17582
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 8342 17370 8402 17582
rect 24577 17579 24643 17582
rect 9949 17506 10015 17509
rect 16389 17506 16455 17509
rect 9949 17504 16455 17506
rect 9949 17448 9954 17504
rect 10010 17448 16394 17504
rect 16450 17448 16455 17504
rect 9949 17446 16455 17448
rect 9949 17443 10015 17446
rect 16389 17443 16455 17446
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 15469 17370 15535 17373
rect 8342 17368 15535 17370
rect 8342 17312 15474 17368
rect 15530 17312 15535 17368
rect 8342 17310 15535 17312
rect 15469 17307 15535 17310
rect 22686 17308 22692 17372
rect 22756 17370 22762 17372
rect 22921 17370 22987 17373
rect 22756 17368 22987 17370
rect 22756 17312 22926 17368
rect 22982 17312 22987 17368
rect 22756 17310 22987 17312
rect 22756 17308 22762 17310
rect 22921 17307 22987 17310
rect 4889 17234 4955 17237
rect 17861 17234 17927 17237
rect 4889 17232 17927 17234
rect 4889 17176 4894 17232
rect 4950 17176 17866 17232
rect 17922 17176 17927 17232
rect 4889 17174 17927 17176
rect 4889 17171 4955 17174
rect 17861 17171 17927 17174
rect 4705 17098 4771 17101
rect 22461 17098 22527 17101
rect 4705 17096 22527 17098
rect 4705 17040 4710 17096
rect 4766 17040 22466 17096
rect 22522 17040 22527 17096
rect 4705 17038 22527 17040
rect 4705 17035 4771 17038
rect 22461 17035 22527 17038
rect 25129 17098 25195 17101
rect 26200 17098 27000 17128
rect 25129 17096 27000 17098
rect 25129 17040 25134 17096
rect 25190 17040 27000 17096
rect 25129 17038 27000 17040
rect 25129 17035 25195 17038
rect 26200 17008 27000 17038
rect 4286 16900 4292 16964
rect 4356 16962 4362 16964
rect 10133 16962 10199 16965
rect 4356 16960 10199 16962
rect 4356 16904 10138 16960
rect 10194 16904 10199 16960
rect 4356 16902 10199 16904
rect 4356 16900 4362 16902
rect 10133 16899 10199 16902
rect 11513 16962 11579 16965
rect 11881 16962 11947 16965
rect 11513 16960 11947 16962
rect 11513 16904 11518 16960
rect 11574 16904 11886 16960
rect 11942 16904 11947 16960
rect 11513 16902 11947 16904
rect 11513 16899 11579 16902
rect 11881 16899 11947 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 7373 16826 7439 16829
rect 7373 16824 12450 16826
rect 7373 16768 7378 16824
rect 7434 16768 12450 16824
rect 7373 16766 12450 16768
rect 7373 16763 7439 16766
rect 6453 16692 6519 16693
rect 8293 16692 8359 16693
rect 9765 16692 9831 16693
rect 6453 16688 6500 16692
rect 6564 16690 6570 16692
rect 8293 16690 8340 16692
rect 6453 16632 6458 16688
rect 6453 16628 6500 16632
rect 6564 16630 6610 16690
rect 8248 16688 8340 16690
rect 8248 16632 8298 16688
rect 8248 16630 8340 16632
rect 6564 16628 6570 16630
rect 8293 16628 8340 16630
rect 8404 16628 8410 16692
rect 9765 16688 9812 16692
rect 9876 16690 9882 16692
rect 12390 16690 12450 16766
rect 16113 16690 16179 16693
rect 9765 16632 9770 16688
rect 9765 16628 9812 16632
rect 9876 16630 9922 16690
rect 12390 16688 16179 16690
rect 12390 16632 16118 16688
rect 16174 16632 16179 16688
rect 12390 16630 16179 16632
rect 9876 16628 9882 16630
rect 6453 16627 6519 16628
rect 8293 16627 8359 16628
rect 9765 16627 9831 16628
rect 16113 16627 16179 16630
rect 16389 16690 16455 16693
rect 17493 16690 17559 16693
rect 16389 16688 17559 16690
rect 16389 16632 16394 16688
rect 16450 16632 17498 16688
rect 17554 16632 17559 16688
rect 16389 16630 17559 16632
rect 16389 16627 16455 16630
rect 17493 16627 17559 16630
rect 7925 16554 7991 16557
rect 18689 16554 18755 16557
rect 7925 16552 18755 16554
rect 7925 16496 7930 16552
rect 7986 16496 18694 16552
rect 18750 16496 18755 16552
rect 7925 16494 18755 16496
rect 7925 16491 7991 16494
rect 18689 16491 18755 16494
rect 8477 16418 8543 16421
rect 9070 16418 9076 16420
rect 8477 16416 9076 16418
rect 8477 16360 8482 16416
rect 8538 16360 9076 16416
rect 8477 16358 9076 16360
rect 8477 16355 8543 16358
rect 9070 16356 9076 16358
rect 9140 16356 9146 16420
rect 11646 16356 11652 16420
rect 11716 16418 11722 16420
rect 12249 16418 12315 16421
rect 11716 16416 12315 16418
rect 11716 16360 12254 16416
rect 12310 16360 12315 16416
rect 11716 16358 12315 16360
rect 11716 16356 11722 16358
rect 12249 16355 12315 16358
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 8886 16220 8892 16284
rect 8956 16282 8962 16284
rect 9029 16282 9095 16285
rect 8956 16280 9095 16282
rect 8956 16224 9034 16280
rect 9090 16224 9095 16280
rect 8956 16222 9095 16224
rect 8956 16220 8962 16222
rect 9029 16219 9095 16222
rect 9949 16282 10015 16285
rect 13997 16282 14063 16285
rect 9949 16280 14063 16282
rect 9949 16224 9954 16280
rect 10010 16224 14002 16280
rect 14058 16224 14063 16280
rect 9949 16222 14063 16224
rect 9949 16219 10015 16222
rect 13997 16219 14063 16222
rect 25037 16282 25103 16285
rect 26200 16282 27000 16312
rect 25037 16280 27000 16282
rect 25037 16224 25042 16280
rect 25098 16224 27000 16280
rect 25037 16222 27000 16224
rect 25037 16219 25103 16222
rect 26200 16192 27000 16222
rect 4981 16146 5047 16149
rect 16665 16146 16731 16149
rect 4981 16144 16731 16146
rect 4981 16088 4986 16144
rect 5042 16088 16670 16144
rect 16726 16088 16731 16144
rect 4981 16086 16731 16088
rect 4981 16083 5047 16086
rect 16665 16083 16731 16086
rect 16849 16146 16915 16149
rect 19742 16146 19748 16148
rect 16849 16144 19748 16146
rect 16849 16088 16854 16144
rect 16910 16088 19748 16144
rect 16849 16086 19748 16088
rect 16849 16083 16915 16086
rect 19742 16084 19748 16086
rect 19812 16084 19818 16148
rect 4061 16010 4127 16013
rect 15285 16010 15351 16013
rect 18505 16010 18571 16013
rect 4061 16008 15210 16010
rect 4061 15952 4066 16008
rect 4122 15952 15210 16008
rect 4061 15950 15210 15952
rect 4061 15947 4127 15950
rect 4429 15874 4495 15877
rect 11237 15874 11303 15877
rect 4429 15872 11303 15874
rect 4429 15816 4434 15872
rect 4490 15816 11242 15872
rect 11298 15816 11303 15872
rect 4429 15814 11303 15816
rect 15150 15874 15210 15950
rect 15285 16008 18571 16010
rect 15285 15952 15290 16008
rect 15346 15952 18510 16008
rect 18566 15952 18571 16008
rect 15285 15950 18571 15952
rect 15285 15947 15351 15950
rect 18505 15947 18571 15950
rect 19374 15874 19380 15876
rect 15150 15814 19380 15874
rect 4429 15811 4495 15814
rect 11237 15811 11303 15814
rect 19374 15812 19380 15814
rect 19444 15812 19450 15876
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 3417 15738 3483 15741
rect 19057 15738 19123 15741
rect 3417 15736 12450 15738
rect 3417 15680 3422 15736
rect 3478 15680 12450 15736
rect 3417 15678 12450 15680
rect 3417 15675 3483 15678
rect 1761 15602 1827 15605
rect 8385 15602 8451 15605
rect 1761 15600 8451 15602
rect 1761 15544 1766 15600
rect 1822 15544 8390 15600
rect 8446 15544 8451 15600
rect 1761 15542 8451 15544
rect 12390 15602 12450 15678
rect 13494 15736 19123 15738
rect 13494 15680 19062 15736
rect 19118 15680 19123 15736
rect 13494 15678 19123 15680
rect 13494 15602 13554 15678
rect 12390 15542 13554 15602
rect 15150 15605 15210 15678
rect 19057 15675 19123 15678
rect 15150 15600 15259 15605
rect 15150 15544 15198 15600
rect 15254 15544 15259 15600
rect 15150 15542 15259 15544
rect 1761 15539 1827 15542
rect 8385 15539 8451 15542
rect 15193 15539 15259 15542
rect 15326 15540 15332 15604
rect 15396 15602 15402 15604
rect 15561 15602 15627 15605
rect 15396 15600 15627 15602
rect 15396 15544 15566 15600
rect 15622 15544 15627 15600
rect 15396 15542 15627 15544
rect 15396 15540 15402 15542
rect 15561 15539 15627 15542
rect 4245 15466 4311 15469
rect 5073 15466 5139 15469
rect 7925 15466 7991 15469
rect 4245 15464 7991 15466
rect 4245 15408 4250 15464
rect 4306 15408 5078 15464
rect 5134 15408 7930 15464
rect 7986 15408 7991 15464
rect 4245 15406 7991 15408
rect 4245 15403 4311 15406
rect 5073 15403 5139 15406
rect 7925 15403 7991 15406
rect 8109 15466 8175 15469
rect 18505 15466 18571 15469
rect 8109 15464 18571 15466
rect 8109 15408 8114 15464
rect 8170 15408 18510 15464
rect 18566 15408 18571 15464
rect 8109 15406 18571 15408
rect 8109 15403 8175 15406
rect 18505 15403 18571 15406
rect 25037 15466 25103 15469
rect 26200 15466 27000 15496
rect 25037 15464 27000 15466
rect 25037 15408 25042 15464
rect 25098 15408 27000 15464
rect 25037 15406 27000 15408
rect 25037 15403 25103 15406
rect 26200 15376 27000 15406
rect 1710 15268 1716 15332
rect 1780 15330 1786 15332
rect 2037 15330 2103 15333
rect 1780 15328 2103 15330
rect 1780 15272 2042 15328
rect 2098 15272 2103 15328
rect 1780 15270 2103 15272
rect 1780 15268 1786 15270
rect 2037 15267 2103 15270
rect 8385 15330 8451 15333
rect 15510 15330 15516 15332
rect 8385 15328 15516 15330
rect 8385 15272 8390 15328
rect 8446 15272 15516 15328
rect 8385 15270 15516 15272
rect 8385 15267 8451 15270
rect 15510 15268 15516 15270
rect 15580 15268 15586 15332
rect 15929 15330 15995 15333
rect 17166 15330 17172 15332
rect 15929 15328 17172 15330
rect 15929 15272 15934 15328
rect 15990 15272 17172 15328
rect 15929 15270 17172 15272
rect 15929 15267 15995 15270
rect 17166 15268 17172 15270
rect 17236 15268 17242 15332
rect 19517 15330 19583 15333
rect 20478 15330 20484 15332
rect 19517 15328 20484 15330
rect 19517 15272 19522 15328
rect 19578 15272 20484 15328
rect 19517 15270 20484 15272
rect 19517 15267 19583 15270
rect 20478 15268 20484 15270
rect 20548 15330 20554 15332
rect 20897 15330 20963 15333
rect 20548 15328 20963 15330
rect 20548 15272 20902 15328
rect 20958 15272 20963 15328
rect 20548 15270 20963 15272
rect 20548 15268 20554 15270
rect 20897 15267 20963 15270
rect 21214 15268 21220 15332
rect 21284 15330 21290 15332
rect 25865 15330 25931 15333
rect 21284 15328 25931 15330
rect 21284 15272 25870 15328
rect 25926 15272 25931 15328
rect 21284 15270 25931 15272
rect 21284 15268 21290 15270
rect 25865 15267 25931 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 7557 15196 7623 15197
rect 7557 15194 7604 15196
rect 7512 15192 7604 15194
rect 7512 15136 7562 15192
rect 7512 15134 7604 15136
rect 7557 15132 7604 15134
rect 7668 15132 7674 15196
rect 10869 15194 10935 15197
rect 14825 15194 14891 15197
rect 10869 15192 14891 15194
rect 10869 15136 10874 15192
rect 10930 15136 14830 15192
rect 14886 15136 14891 15192
rect 10869 15134 14891 15136
rect 7557 15131 7623 15132
rect 10869 15131 10935 15134
rect 14825 15131 14891 15134
rect 24669 15196 24735 15197
rect 24669 15192 24716 15196
rect 24780 15194 24786 15196
rect 24669 15136 24674 15192
rect 24669 15132 24716 15136
rect 24780 15134 24826 15194
rect 24780 15132 24786 15134
rect 24669 15131 24735 15132
rect 7189 15058 7255 15061
rect 7925 15058 7991 15061
rect 7189 15056 7991 15058
rect 7189 15000 7194 15056
rect 7250 15000 7930 15056
rect 7986 15000 7991 15056
rect 7189 14998 7991 15000
rect 7189 14995 7255 14998
rect 7925 14995 7991 14998
rect 12750 14996 12756 15060
rect 12820 15058 12826 15060
rect 20345 15058 20411 15061
rect 12820 15056 20411 15058
rect 12820 15000 20350 15056
rect 20406 15000 20411 15056
rect 12820 14998 20411 15000
rect 12820 14996 12826 14998
rect 20345 14995 20411 14998
rect 1158 14860 1164 14924
rect 1228 14922 1234 14924
rect 3233 14922 3299 14925
rect 1228 14920 3299 14922
rect 1228 14864 3238 14920
rect 3294 14864 3299 14920
rect 1228 14862 3299 14864
rect 1228 14860 1234 14862
rect 3233 14859 3299 14862
rect 6545 14922 6611 14925
rect 21633 14922 21699 14925
rect 6545 14920 21699 14922
rect 6545 14864 6550 14920
rect 6606 14864 21638 14920
rect 21694 14864 21699 14920
rect 6545 14862 21699 14864
rect 6545 14859 6611 14862
rect 21633 14859 21699 14862
rect 3785 14786 3851 14789
rect 11329 14786 11395 14789
rect 3785 14784 11395 14786
rect 3785 14728 3790 14784
rect 3846 14728 11334 14784
rect 11390 14728 11395 14784
rect 3785 14726 11395 14728
rect 3785 14723 3851 14726
rect 11329 14723 11395 14726
rect 17534 14724 17540 14788
rect 17604 14786 17610 14788
rect 19793 14786 19859 14789
rect 17604 14784 19859 14786
rect 17604 14728 19798 14784
rect 19854 14728 19859 14784
rect 17604 14726 19859 14728
rect 17604 14724 17610 14726
rect 19793 14723 19859 14726
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 6545 14650 6611 14653
rect 12750 14650 12756 14652
rect 6545 14648 12756 14650
rect 6545 14592 6550 14648
rect 6606 14592 12756 14648
rect 6545 14590 12756 14592
rect 6545 14587 6611 14590
rect 12750 14588 12756 14590
rect 12820 14588 12826 14652
rect 21725 14650 21791 14653
rect 22134 14650 22140 14652
rect 21725 14648 22140 14650
rect 21725 14592 21730 14648
rect 21786 14592 22140 14648
rect 21725 14590 22140 14592
rect 21725 14587 21791 14590
rect 22134 14588 22140 14590
rect 22204 14588 22210 14652
rect 23381 14650 23447 14653
rect 26200 14650 27000 14680
rect 23381 14648 27000 14650
rect 23381 14592 23386 14648
rect 23442 14592 27000 14648
rect 23381 14590 27000 14592
rect 23381 14587 23447 14590
rect 26200 14560 27000 14590
rect 6269 14514 6335 14517
rect 6269 14512 22064 14514
rect 6269 14456 6274 14512
rect 6330 14456 22064 14512
rect 6269 14454 22064 14456
rect 6269 14451 6335 14454
rect 22004 14381 22064 14454
rect 5257 14378 5323 14381
rect 21265 14378 21331 14381
rect 5257 14376 21331 14378
rect 5257 14320 5262 14376
rect 5318 14320 21270 14376
rect 21326 14320 21331 14376
rect 5257 14318 21331 14320
rect 5257 14315 5323 14318
rect 21265 14315 21331 14318
rect 22001 14376 22067 14381
rect 22001 14320 22006 14376
rect 22062 14320 22067 14376
rect 22001 14315 22067 14320
rect 2037 14242 2103 14245
rect 5574 14242 5580 14244
rect 2037 14240 5580 14242
rect 2037 14184 2042 14240
rect 2098 14184 5580 14240
rect 2037 14182 5580 14184
rect 2037 14179 2103 14182
rect 5574 14180 5580 14182
rect 5644 14180 5650 14244
rect 11237 14242 11303 14245
rect 16389 14244 16455 14245
rect 13854 14242 13860 14244
rect 11237 14240 13860 14242
rect 11237 14184 11242 14240
rect 11298 14184 13860 14240
rect 11237 14182 13860 14184
rect 11237 14179 11303 14182
rect 13854 14180 13860 14182
rect 13924 14180 13930 14244
rect 16389 14242 16436 14244
rect 16344 14240 16436 14242
rect 16344 14184 16394 14240
rect 16344 14182 16436 14184
rect 16389 14180 16436 14182
rect 16500 14180 16506 14244
rect 16614 14180 16620 14244
rect 16684 14242 16690 14244
rect 16849 14242 16915 14245
rect 16684 14240 16915 14242
rect 16684 14184 16854 14240
rect 16910 14184 16915 14240
rect 16684 14182 16915 14184
rect 16684 14180 16690 14182
rect 16389 14179 16455 14180
rect 16849 14179 16915 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 10869 14106 10935 14109
rect 12566 14106 12572 14108
rect 10869 14104 12572 14106
rect 10869 14048 10874 14104
rect 10930 14048 12572 14104
rect 10869 14046 12572 14048
rect 10869 14043 10935 14046
rect 12566 14044 12572 14046
rect 12636 14044 12642 14108
rect 16481 14106 16547 14109
rect 13494 14104 16547 14106
rect 13494 14048 16486 14104
rect 16542 14048 16547 14104
rect 13494 14046 16547 14048
rect 1853 13970 1919 13973
rect 3785 13970 3851 13973
rect 1853 13968 3851 13970
rect 1853 13912 1858 13968
rect 1914 13912 3790 13968
rect 3846 13912 3851 13968
rect 1853 13910 3851 13912
rect 1853 13907 1919 13910
rect 3785 13907 3851 13910
rect 4061 13970 4127 13973
rect 13494 13970 13554 14046
rect 16481 14043 16547 14046
rect 4061 13968 13554 13970
rect 4061 13912 4066 13968
rect 4122 13912 13554 13968
rect 4061 13910 13554 13912
rect 4061 13907 4127 13910
rect 13670 13908 13676 13972
rect 13740 13970 13746 13972
rect 20437 13970 20503 13973
rect 13740 13968 20503 13970
rect 13740 13912 20442 13968
rect 20498 13912 20503 13968
rect 13740 13910 20503 13912
rect 13740 13908 13746 13910
rect 20437 13907 20503 13910
rect 2446 13772 2452 13836
rect 2516 13834 2522 13836
rect 2589 13834 2655 13837
rect 2516 13832 2655 13834
rect 2516 13776 2594 13832
rect 2650 13776 2655 13832
rect 2516 13774 2655 13776
rect 2516 13772 2522 13774
rect 2589 13771 2655 13774
rect 6913 13834 6979 13837
rect 15193 13834 15259 13837
rect 6913 13832 15259 13834
rect 6913 13776 6918 13832
rect 6974 13776 15198 13832
rect 15254 13776 15259 13832
rect 6913 13774 15259 13776
rect 6913 13771 6979 13774
rect 15193 13771 15259 13774
rect 16481 13834 16547 13837
rect 20662 13834 20668 13836
rect 16481 13832 20668 13834
rect 16481 13776 16486 13832
rect 16542 13776 20668 13832
rect 16481 13774 20668 13776
rect 16481 13771 16547 13774
rect 20662 13772 20668 13774
rect 20732 13772 20738 13836
rect 23933 13834 23999 13837
rect 26200 13834 27000 13864
rect 23933 13832 27000 13834
rect 23933 13776 23938 13832
rect 23994 13776 27000 13832
rect 23933 13774 27000 13776
rect 23933 13771 23999 13774
rect 26200 13744 27000 13774
rect 3417 13700 3483 13701
rect 3366 13636 3372 13700
rect 3436 13698 3483 13700
rect 13353 13698 13419 13701
rect 16113 13698 16179 13701
rect 17769 13700 17835 13701
rect 17718 13698 17724 13700
rect 3436 13696 12450 13698
rect 3478 13640 12450 13696
rect 3436 13638 12450 13640
rect 3436 13636 3483 13638
rect 3417 13635 3483 13636
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 5758 13500 5764 13564
rect 5828 13562 5834 13564
rect 9949 13562 10015 13565
rect 12390 13564 12450 13638
rect 13353 13696 16179 13698
rect 13353 13640 13358 13696
rect 13414 13640 16118 13696
rect 16174 13640 16179 13696
rect 13353 13638 16179 13640
rect 17678 13638 17724 13698
rect 17788 13696 17835 13700
rect 17830 13640 17835 13696
rect 13353 13635 13419 13638
rect 16113 13635 16179 13638
rect 17718 13636 17724 13638
rect 17788 13636 17835 13640
rect 17769 13635 17835 13636
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 5828 13560 10015 13562
rect 5828 13504 9954 13560
rect 10010 13504 10015 13560
rect 5828 13502 10015 13504
rect 5828 13500 5834 13502
rect 9949 13499 10015 13502
rect 12382 13500 12388 13564
rect 12452 13500 12458 13564
rect 15469 13562 15535 13565
rect 15837 13562 15903 13565
rect 19333 13564 19399 13565
rect 19333 13562 19380 13564
rect 15469 13560 15903 13562
rect 15469 13504 15474 13560
rect 15530 13504 15842 13560
rect 15898 13504 15903 13560
rect 15469 13502 15903 13504
rect 19288 13560 19380 13562
rect 19288 13504 19338 13560
rect 19288 13502 19380 13504
rect 15469 13499 15535 13502
rect 15837 13499 15903 13502
rect 19333 13500 19380 13502
rect 19444 13500 19450 13564
rect 19333 13499 19399 13500
rect 4245 13426 4311 13429
rect 20621 13426 20687 13429
rect 4245 13424 20687 13426
rect 4245 13368 4250 13424
rect 4306 13368 20626 13424
rect 20682 13368 20687 13424
rect 4245 13366 20687 13368
rect 4245 13363 4311 13366
rect 20621 13363 20687 13366
rect 5165 13290 5231 13293
rect 12065 13290 12131 13293
rect 12198 13290 12204 13292
rect 5165 13288 8770 13290
rect 5165 13232 5170 13288
rect 5226 13232 8770 13288
rect 5165 13230 8770 13232
rect 5165 13227 5231 13230
rect 8710 13154 8770 13230
rect 12065 13288 12204 13290
rect 12065 13232 12070 13288
rect 12126 13232 12204 13288
rect 12065 13230 12204 13232
rect 12065 13227 12131 13230
rect 12198 13228 12204 13230
rect 12268 13228 12274 13292
rect 12382 13228 12388 13292
rect 12452 13290 12458 13292
rect 20713 13290 20779 13293
rect 24577 13292 24643 13293
rect 12452 13288 20779 13290
rect 12452 13232 20718 13288
rect 20774 13232 20779 13288
rect 12452 13230 20779 13232
rect 12452 13228 12458 13230
rect 20713 13227 20779 13230
rect 24526 13228 24532 13292
rect 24596 13290 24643 13292
rect 24596 13288 24688 13290
rect 24638 13232 24688 13288
rect 24596 13230 24688 13232
rect 24596 13228 24643 13230
rect 24577 13227 24643 13228
rect 8710 13094 17280 13154
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 9765 13018 9831 13021
rect 11697 13018 11763 13021
rect 9765 13016 11763 13018
rect 9765 12960 9770 13016
rect 9826 12960 11702 13016
rect 11758 12960 11763 13016
rect 9765 12958 11763 12960
rect 9765 12955 9831 12958
rect 11697 12955 11763 12958
rect 12341 13018 12407 13021
rect 15469 13018 15535 13021
rect 16113 13018 16179 13021
rect 12341 13016 16179 13018
rect 12341 12960 12346 13016
rect 12402 12960 15474 13016
rect 15530 12960 16118 13016
rect 16174 12960 16179 13016
rect 12341 12958 16179 12960
rect 12341 12955 12407 12958
rect 15469 12955 15535 12958
rect 16113 12955 16179 12958
rect 5073 12882 5139 12885
rect 17220 12882 17280 13094
rect 19190 13092 19196 13156
rect 19260 13154 19266 13156
rect 19517 13154 19583 13157
rect 19260 13152 19583 13154
rect 19260 13096 19522 13152
rect 19578 13096 19583 13152
rect 19260 13094 19583 13096
rect 19260 13092 19266 13094
rect 19517 13091 19583 13094
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 22093 13020 22159 13021
rect 22093 13018 22140 13020
rect 22048 13016 22140 13018
rect 22048 12960 22098 13016
rect 22048 12958 22140 12960
rect 22093 12956 22140 12958
rect 22204 12956 22210 13020
rect 24761 13018 24827 13021
rect 26200 13018 27000 13048
rect 24761 13016 27000 13018
rect 24761 12960 24766 13016
rect 24822 12960 27000 13016
rect 24761 12958 27000 12960
rect 22093 12955 22159 12956
rect 24761 12955 24827 12958
rect 26200 12928 27000 12958
rect 23289 12882 23355 12885
rect 23933 12882 23999 12885
rect 5073 12880 17050 12882
rect 5073 12824 5078 12880
rect 5134 12824 17050 12880
rect 5073 12822 17050 12824
rect 17220 12880 23999 12882
rect 17220 12824 23294 12880
rect 23350 12824 23938 12880
rect 23994 12824 23999 12880
rect 17220 12822 23999 12824
rect 5073 12819 5139 12822
rect 1761 12746 1827 12749
rect 4470 12746 4476 12748
rect 1761 12744 4476 12746
rect 1761 12688 1766 12744
rect 1822 12688 4476 12744
rect 1761 12686 4476 12688
rect 1761 12683 1827 12686
rect 4470 12684 4476 12686
rect 4540 12684 4546 12748
rect 5533 12746 5599 12749
rect 16990 12746 17050 12822
rect 23289 12819 23355 12822
rect 23933 12819 23999 12822
rect 21449 12746 21515 12749
rect 5533 12744 16636 12746
rect 5533 12688 5538 12744
rect 5594 12688 16636 12744
rect 5533 12686 16636 12688
rect 16990 12744 21515 12746
rect 16990 12688 21454 12744
rect 21510 12688 21515 12744
rect 16990 12686 21515 12688
rect 5533 12683 5599 12686
rect 3785 12610 3851 12613
rect 3918 12610 3924 12612
rect 3785 12608 3924 12610
rect 3785 12552 3790 12608
rect 3846 12552 3924 12608
rect 3785 12550 3924 12552
rect 3785 12547 3851 12550
rect 3918 12548 3924 12550
rect 3988 12548 3994 12612
rect 5625 12610 5691 12613
rect 6177 12610 6243 12613
rect 5625 12608 6243 12610
rect 5625 12552 5630 12608
rect 5686 12552 6182 12608
rect 6238 12552 6243 12608
rect 5625 12550 6243 12552
rect 5625 12547 5691 12550
rect 6177 12547 6243 12550
rect 6637 12610 6703 12613
rect 13721 12610 13787 12613
rect 15561 12610 15627 12613
rect 6637 12608 12818 12610
rect 6637 12552 6642 12608
rect 6698 12552 12818 12608
rect 6637 12550 12818 12552
rect 6637 12547 6703 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 3601 12474 3667 12477
rect 7557 12474 7623 12477
rect 3601 12472 7623 12474
rect 3601 12416 3606 12472
rect 3662 12416 7562 12472
rect 7618 12416 7623 12472
rect 3601 12414 7623 12416
rect 3601 12411 3667 12414
rect 7557 12411 7623 12414
rect 8753 12474 8819 12477
rect 10133 12474 10199 12477
rect 8753 12472 10199 12474
rect 8753 12416 8758 12472
rect 8814 12416 10138 12472
rect 10194 12416 10199 12472
rect 8753 12414 10199 12416
rect 8753 12411 8819 12414
rect 10133 12411 10199 12414
rect 11697 12474 11763 12477
rect 12157 12474 12223 12477
rect 11697 12472 12223 12474
rect 11697 12416 11702 12472
rect 11758 12416 12162 12472
rect 12218 12416 12223 12472
rect 11697 12414 12223 12416
rect 11697 12411 11763 12414
rect 12157 12411 12223 12414
rect 2129 12340 2195 12341
rect 2078 12276 2084 12340
rect 2148 12338 2195 12340
rect 4061 12338 4127 12341
rect 11605 12338 11671 12341
rect 2148 12336 2240 12338
rect 2190 12280 2240 12336
rect 2148 12278 2240 12280
rect 4061 12336 11671 12338
rect 4061 12280 4066 12336
rect 4122 12280 11610 12336
rect 11666 12280 11671 12336
rect 4061 12278 11671 12280
rect 12758 12338 12818 12550
rect 13721 12608 15627 12610
rect 13721 12552 13726 12608
rect 13782 12552 15566 12608
rect 15622 12552 15627 12608
rect 13721 12550 15627 12552
rect 13721 12547 13787 12550
rect 15561 12547 15627 12550
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 16389 12474 16455 12477
rect 13356 12472 16455 12474
rect 13356 12416 16394 12472
rect 16450 12416 16455 12472
rect 13356 12414 16455 12416
rect 16576 12474 16636 12686
rect 21449 12683 21515 12686
rect 20713 12610 20779 12613
rect 21214 12610 21220 12612
rect 20713 12608 21220 12610
rect 20713 12552 20718 12608
rect 20774 12552 21220 12608
rect 20713 12550 21220 12552
rect 20713 12547 20779 12550
rect 21214 12548 21220 12550
rect 21284 12548 21290 12612
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 18321 12474 18387 12477
rect 20989 12474 21055 12477
rect 16576 12472 21055 12474
rect 16576 12416 18326 12472
rect 18382 12416 20994 12472
rect 21050 12416 21055 12472
rect 16576 12414 21055 12416
rect 13356 12338 13416 12414
rect 16389 12411 16455 12414
rect 18321 12411 18387 12414
rect 20989 12411 21055 12414
rect 12758 12278 13416 12338
rect 13629 12338 13695 12341
rect 17493 12338 17559 12341
rect 13629 12336 17559 12338
rect 13629 12280 13634 12336
rect 13690 12280 17498 12336
rect 17554 12280 17559 12336
rect 13629 12278 17559 12280
rect 2148 12276 2195 12278
rect 2129 12275 2195 12276
rect 4061 12275 4127 12278
rect 11605 12275 11671 12278
rect 13629 12275 13695 12278
rect 17493 12275 17559 12278
rect 2129 12202 2195 12205
rect 16481 12202 16547 12205
rect 2129 12200 16547 12202
rect 2129 12144 2134 12200
rect 2190 12144 16486 12200
rect 16542 12144 16547 12200
rect 2129 12142 16547 12144
rect 2129 12139 2195 12142
rect 16481 12139 16547 12142
rect 24853 12202 24919 12205
rect 26200 12202 27000 12232
rect 24853 12200 27000 12202
rect 24853 12144 24858 12200
rect 24914 12144 27000 12200
rect 24853 12142 27000 12144
rect 24853 12139 24919 12142
rect 26200 12112 27000 12142
rect 9673 12066 9739 12069
rect 14917 12066 14983 12069
rect 9673 12064 14983 12066
rect 9673 12008 9678 12064
rect 9734 12008 14922 12064
rect 14978 12008 14983 12064
rect 9673 12006 14983 12008
rect 9673 12003 9739 12006
rect 14917 12003 14983 12006
rect 16573 12066 16639 12069
rect 17677 12066 17743 12069
rect 16573 12064 17743 12066
rect 16573 12008 16578 12064
rect 16634 12008 17682 12064
rect 17738 12008 17743 12064
rect 16573 12006 17743 12008
rect 16573 12003 16639 12006
rect 17677 12003 17743 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 10501 11930 10567 11933
rect 11973 11930 12039 11933
rect 10501 11928 12039 11930
rect 10501 11872 10506 11928
rect 10562 11872 11978 11928
rect 12034 11872 12039 11928
rect 10501 11870 12039 11872
rect 10501 11867 10567 11870
rect 11973 11867 12039 11870
rect 12750 11868 12756 11932
rect 12820 11930 12826 11932
rect 15694 11930 15700 11932
rect 12820 11870 15700 11930
rect 12820 11868 12826 11870
rect 15694 11868 15700 11870
rect 15764 11868 15770 11932
rect 3969 11794 4035 11797
rect 17217 11794 17283 11797
rect 3969 11792 17283 11794
rect 3969 11736 3974 11792
rect 4030 11736 17222 11792
rect 17278 11736 17283 11792
rect 3969 11734 17283 11736
rect 3969 11731 4035 11734
rect 17217 11731 17283 11734
rect 20662 11732 20668 11796
rect 20732 11794 20738 11796
rect 23749 11794 23815 11797
rect 20732 11792 23815 11794
rect 20732 11736 23754 11792
rect 23810 11736 23815 11792
rect 20732 11734 23815 11736
rect 20732 11732 20738 11734
rect 23749 11731 23815 11734
rect 5993 11658 6059 11661
rect 23289 11658 23355 11661
rect 5993 11656 23355 11658
rect 5993 11600 5998 11656
rect 6054 11600 23294 11656
rect 23350 11600 23355 11656
rect 5993 11598 23355 11600
rect 5993 11595 6059 11598
rect 23289 11595 23355 11598
rect 6913 11522 6979 11525
rect 8334 11522 8340 11524
rect 6913 11520 8340 11522
rect 6913 11464 6918 11520
rect 6974 11464 8340 11520
rect 6913 11462 8340 11464
rect 6913 11459 6979 11462
rect 8334 11460 8340 11462
rect 8404 11460 8410 11524
rect 10317 11522 10383 11525
rect 12709 11522 12775 11525
rect 10317 11520 12775 11522
rect 10317 11464 10322 11520
rect 10378 11464 12714 11520
rect 12770 11464 12775 11520
rect 10317 11462 12775 11464
rect 10317 11459 10383 11462
rect 12709 11459 12775 11462
rect 15326 11460 15332 11524
rect 15396 11522 15402 11524
rect 19701 11522 19767 11525
rect 15396 11520 19767 11522
rect 15396 11464 19706 11520
rect 19762 11464 19767 11520
rect 15396 11462 19767 11464
rect 15396 11460 15402 11462
rect 19701 11459 19767 11462
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 8293 11386 8359 11389
rect 12750 11386 12756 11388
rect 8293 11384 12756 11386
rect 8293 11328 8298 11384
rect 8354 11328 12756 11384
rect 8293 11326 12756 11328
rect 8293 11323 8359 11326
rect 12750 11324 12756 11326
rect 12820 11324 12826 11388
rect 13629 11386 13695 11389
rect 17861 11386 17927 11389
rect 13629 11384 17927 11386
rect 13629 11328 13634 11384
rect 13690 11328 17866 11384
rect 17922 11328 17927 11384
rect 13629 11326 17927 11328
rect 13629 11323 13695 11326
rect 17861 11323 17927 11326
rect 19333 11386 19399 11389
rect 19742 11386 19748 11388
rect 19333 11384 19748 11386
rect 19333 11328 19338 11384
rect 19394 11328 19748 11384
rect 19333 11326 19748 11328
rect 19333 11323 19399 11326
rect 19742 11324 19748 11326
rect 19812 11324 19818 11388
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 7465 11250 7531 11253
rect 16573 11250 16639 11253
rect 18965 11250 19031 11253
rect 7465 11248 16639 11250
rect 7465 11192 7470 11248
rect 7526 11192 16578 11248
rect 16634 11192 16639 11248
rect 7465 11190 16639 11192
rect 7465 11187 7531 11190
rect 16573 11187 16639 11190
rect 17358 11248 19031 11250
rect 17358 11192 18970 11248
rect 19026 11192 19031 11248
rect 17358 11190 19031 11192
rect 3233 11114 3299 11117
rect 17358 11114 17418 11190
rect 18965 11187 19031 11190
rect 20161 11250 20227 11253
rect 23657 11250 23723 11253
rect 20161 11248 23723 11250
rect 20161 11192 20166 11248
rect 20222 11192 23662 11248
rect 23718 11192 23723 11248
rect 20161 11190 23723 11192
rect 20161 11187 20227 11190
rect 23657 11187 23723 11190
rect 3233 11112 17418 11114
rect 3233 11056 3238 11112
rect 3294 11056 17418 11112
rect 3233 11054 17418 11056
rect 18689 11114 18755 11117
rect 19006 11114 19012 11116
rect 18689 11112 19012 11114
rect 18689 11056 18694 11112
rect 18750 11056 19012 11112
rect 18689 11054 19012 11056
rect 3233 11051 3299 11054
rect 18689 11051 18755 11054
rect 19006 11052 19012 11054
rect 19076 11052 19082 11116
rect 21030 11052 21036 11116
rect 21100 11114 21106 11116
rect 21633 11114 21699 11117
rect 21100 11112 21699 11114
rect 21100 11056 21638 11112
rect 21694 11056 21699 11112
rect 21100 11054 21699 11056
rect 21100 11052 21106 11054
rect 21633 11051 21699 11054
rect 2037 10978 2103 10981
rect 16297 10978 16363 10981
rect 2037 10976 3434 10978
rect 2037 10920 2042 10976
rect 2098 10920 3434 10976
rect 2037 10918 3434 10920
rect 2037 10915 2103 10918
rect 3374 10434 3434 10918
rect 8342 10976 16363 10978
rect 8342 10920 16302 10976
rect 16358 10920 16363 10976
rect 8342 10918 16363 10920
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 7281 10706 7347 10709
rect 8342 10706 8402 10918
rect 16297 10915 16363 10918
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 10593 10842 10659 10845
rect 13486 10842 13492 10844
rect 10593 10840 13492 10842
rect 10593 10784 10598 10840
rect 10654 10784 13492 10840
rect 10593 10782 13492 10784
rect 10593 10779 10659 10782
rect 13486 10780 13492 10782
rect 13556 10780 13562 10844
rect 7281 10704 8402 10706
rect 7281 10648 7286 10704
rect 7342 10648 8402 10704
rect 7281 10646 8402 10648
rect 8477 10706 8543 10709
rect 19149 10706 19215 10709
rect 8477 10704 19215 10706
rect 8477 10648 8482 10704
rect 8538 10648 19154 10704
rect 19210 10648 19215 10704
rect 8477 10646 19215 10648
rect 7281 10643 7347 10646
rect 8477 10643 8543 10646
rect 19149 10643 19215 10646
rect 3601 10570 3667 10573
rect 22737 10570 22803 10573
rect 3601 10568 22803 10570
rect 3601 10512 3606 10568
rect 3662 10512 22742 10568
rect 22798 10512 22803 10568
rect 3601 10510 22803 10512
rect 3601 10507 3667 10510
rect 22737 10507 22803 10510
rect 24761 10570 24827 10573
rect 26200 10570 27000 10600
rect 24761 10568 27000 10570
rect 24761 10512 24766 10568
rect 24822 10512 27000 10568
rect 24761 10510 27000 10512
rect 24761 10507 24827 10510
rect 26200 10480 27000 10510
rect 3601 10434 3667 10437
rect 11421 10434 11487 10437
rect 3374 10432 3667 10434
rect 3374 10376 3606 10432
rect 3662 10376 3667 10432
rect 3374 10374 3667 10376
rect 3601 10371 3667 10374
rect 3788 10432 11487 10434
rect 3788 10376 11426 10432
rect 11482 10376 11487 10432
rect 3788 10374 11487 10376
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 2681 10162 2747 10165
rect 3788 10162 3848 10374
rect 11421 10371 11487 10374
rect 11789 10434 11855 10437
rect 12709 10434 12775 10437
rect 11789 10432 12775 10434
rect 11789 10376 11794 10432
rect 11850 10376 12714 10432
rect 12770 10376 12775 10432
rect 11789 10374 12775 10376
rect 11789 10371 11855 10374
rect 12709 10371 12775 10374
rect 14222 10372 14228 10436
rect 14292 10434 14298 10436
rect 19190 10434 19196 10436
rect 14292 10374 19196 10434
rect 14292 10372 14298 10374
rect 19190 10372 19196 10374
rect 19260 10372 19266 10436
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 4245 10298 4311 10301
rect 7005 10298 7071 10301
rect 4245 10296 7071 10298
rect 4245 10240 4250 10296
rect 4306 10240 7010 10296
rect 7066 10240 7071 10296
rect 4245 10238 7071 10240
rect 4245 10235 4311 10238
rect 7005 10235 7071 10238
rect 7230 10236 7236 10300
rect 7300 10298 7306 10300
rect 11094 10298 11100 10300
rect 7300 10238 11100 10298
rect 7300 10236 7306 10238
rect 11094 10236 11100 10238
rect 11164 10236 11170 10300
rect 11605 10298 11671 10301
rect 12750 10298 12756 10300
rect 11605 10296 12756 10298
rect 11605 10240 11610 10296
rect 11666 10240 12756 10296
rect 11605 10238 12756 10240
rect 11605 10235 11671 10238
rect 12750 10236 12756 10238
rect 12820 10236 12826 10300
rect 14457 10298 14523 10301
rect 14917 10298 14983 10301
rect 14457 10296 14983 10298
rect 14457 10240 14462 10296
rect 14518 10240 14922 10296
rect 14978 10240 14983 10296
rect 14457 10238 14983 10240
rect 14457 10235 14523 10238
rect 14917 10235 14983 10238
rect 2681 10160 3848 10162
rect 2681 10104 2686 10160
rect 2742 10104 3848 10160
rect 2681 10102 3848 10104
rect 6637 10162 6703 10165
rect 17861 10162 17927 10165
rect 6637 10160 17927 10162
rect 6637 10104 6642 10160
rect 6698 10104 17866 10160
rect 17922 10104 17927 10160
rect 6637 10102 17927 10104
rect 2681 10099 2747 10102
rect 6637 10099 6703 10102
rect 17861 10099 17927 10102
rect 3233 10026 3299 10029
rect 23197 10026 23263 10029
rect 3233 10024 23263 10026
rect 3233 9968 3238 10024
rect 3294 9968 23202 10024
rect 23258 9968 23263 10024
rect 3233 9966 23263 9968
rect 3233 9963 3299 9966
rect 23197 9963 23263 9966
rect 2681 9890 2747 9893
rect 3366 9890 3372 9892
rect 2681 9888 3372 9890
rect 2681 9832 2686 9888
rect 2742 9832 3372 9888
rect 2681 9830 3372 9832
rect 2681 9827 2747 9830
rect 3366 9828 3372 9830
rect 3436 9828 3442 9892
rect 4981 9890 5047 9893
rect 7230 9890 7236 9892
rect 4981 9888 7236 9890
rect 4981 9832 4986 9888
rect 5042 9832 7236 9888
rect 4981 9830 7236 9832
rect 4981 9827 5047 9830
rect 7230 9828 7236 9830
rect 7300 9828 7306 9892
rect 9581 9890 9647 9893
rect 16389 9890 16455 9893
rect 9581 9888 16455 9890
rect 9581 9832 9586 9888
rect 9642 9832 16394 9888
rect 16450 9832 16455 9888
rect 9581 9830 16455 9832
rect 9581 9827 9647 9830
rect 16389 9827 16455 9830
rect 20253 9890 20319 9893
rect 23841 9890 23907 9893
rect 20253 9888 23907 9890
rect 20253 9832 20258 9888
rect 20314 9832 23846 9888
rect 23902 9832 23907 9888
rect 20253 9830 23907 9832
rect 20253 9827 20319 9830
rect 23841 9827 23907 9830
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 974 9692 980 9756
rect 1044 9754 1050 9756
rect 2037 9754 2103 9757
rect 1044 9752 2103 9754
rect 1044 9696 2042 9752
rect 2098 9696 2103 9752
rect 1044 9694 2103 9696
rect 1044 9692 1050 9694
rect 2037 9691 2103 9694
rect 10409 9754 10475 9757
rect 13169 9754 13235 9757
rect 10409 9752 13235 9754
rect 10409 9696 10414 9752
rect 10470 9696 13174 9752
rect 13230 9696 13235 9752
rect 10409 9694 13235 9696
rect 10409 9691 10475 9694
rect 13169 9691 13235 9694
rect 13813 9754 13879 9757
rect 16614 9754 16620 9756
rect 13813 9752 16620 9754
rect 13813 9696 13818 9752
rect 13874 9696 16620 9752
rect 13813 9694 16620 9696
rect 13813 9691 13879 9694
rect 16614 9692 16620 9694
rect 16684 9692 16690 9756
rect 25129 9754 25195 9757
rect 26200 9754 27000 9784
rect 16806 9694 17234 9754
rect 3233 9618 3299 9621
rect 16806 9618 16866 9694
rect 3233 9616 16866 9618
rect 3233 9560 3238 9616
rect 3294 9560 16866 9616
rect 3233 9558 16866 9560
rect 16941 9620 17007 9621
rect 16941 9616 16988 9620
rect 17052 9618 17058 9620
rect 17174 9618 17234 9694
rect 25129 9752 27000 9754
rect 25129 9696 25134 9752
rect 25190 9696 27000 9752
rect 25129 9694 27000 9696
rect 25129 9691 25195 9694
rect 26200 9664 27000 9694
rect 21081 9618 21147 9621
rect 21725 9618 21791 9621
rect 16941 9560 16946 9616
rect 3233 9555 3299 9558
rect 16941 9556 16988 9560
rect 17052 9558 17098 9618
rect 17174 9616 21791 9618
rect 17174 9560 21086 9616
rect 21142 9560 21730 9616
rect 21786 9560 21791 9616
rect 17174 9558 21791 9560
rect 17052 9556 17058 9558
rect 16941 9555 17007 9556
rect 21081 9555 21147 9558
rect 21725 9555 21791 9558
rect 1853 9482 1919 9485
rect 3366 9482 3372 9484
rect 1853 9480 3372 9482
rect 1853 9424 1858 9480
rect 1914 9424 3372 9480
rect 1853 9422 3372 9424
rect 1853 9419 1919 9422
rect 3366 9420 3372 9422
rect 3436 9482 3442 9484
rect 19977 9482 20043 9485
rect 3436 9480 20043 9482
rect 3436 9424 19982 9480
rect 20038 9424 20043 9480
rect 3436 9422 20043 9424
rect 3436 9420 3442 9422
rect 19977 9419 20043 9422
rect 8201 9346 8267 9349
rect 8518 9346 8524 9348
rect 8201 9344 8524 9346
rect 8201 9288 8206 9344
rect 8262 9288 8524 9344
rect 8201 9286 8524 9288
rect 8201 9283 8267 9286
rect 8518 9284 8524 9286
rect 8588 9284 8594 9348
rect 13854 9284 13860 9348
rect 13924 9346 13930 9348
rect 14181 9346 14247 9349
rect 14365 9346 14431 9349
rect 13924 9344 14431 9346
rect 13924 9288 14186 9344
rect 14242 9288 14370 9344
rect 14426 9288 14431 9344
rect 13924 9286 14431 9288
rect 13924 9284 13930 9286
rect 14181 9283 14247 9286
rect 14365 9283 14431 9286
rect 14590 9284 14596 9348
rect 14660 9346 14666 9348
rect 16021 9346 16087 9349
rect 14660 9344 16087 9346
rect 14660 9288 16026 9344
rect 16082 9288 16087 9344
rect 14660 9286 16087 9288
rect 14660 9284 14666 9286
rect 16021 9283 16087 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 5574 9148 5580 9212
rect 5644 9210 5650 9212
rect 8477 9210 8543 9213
rect 5644 9208 8543 9210
rect 5644 9152 8482 9208
rect 8538 9152 8543 9208
rect 5644 9150 8543 9152
rect 5644 9148 5650 9150
rect 8477 9147 8543 9150
rect 3417 9074 3483 9077
rect 5758 9074 5764 9076
rect 3417 9072 5764 9074
rect 3417 9016 3422 9072
rect 3478 9016 5764 9072
rect 3417 9014 5764 9016
rect 3417 9011 3483 9014
rect 5758 9012 5764 9014
rect 5828 9012 5834 9076
rect 8845 9074 8911 9077
rect 18689 9074 18755 9077
rect 5950 9014 8586 9074
rect 3969 8938 4035 8941
rect 4102 8938 4108 8940
rect 3969 8936 4108 8938
rect 3969 8880 3974 8936
rect 4030 8880 4108 8936
rect 3969 8878 4108 8880
rect 3969 8875 4035 8878
rect 4102 8876 4108 8878
rect 4172 8876 4178 8940
rect 5441 8938 5507 8941
rect 5950 8938 6010 9014
rect 5441 8936 6010 8938
rect 5441 8880 5446 8936
rect 5502 8880 6010 8936
rect 5441 8878 6010 8880
rect 6821 8938 6887 8941
rect 8526 8938 8586 9014
rect 8845 9072 18755 9074
rect 8845 9016 8850 9072
rect 8906 9016 18694 9072
rect 18750 9016 18755 9072
rect 8845 9014 18755 9016
rect 8845 9011 8911 9014
rect 18689 9011 18755 9014
rect 22093 8938 22159 8941
rect 6821 8936 8402 8938
rect 6821 8880 6826 8936
rect 6882 8880 8402 8936
rect 6821 8878 8402 8880
rect 8526 8936 22159 8938
rect 8526 8880 22098 8936
rect 22154 8880 22159 8936
rect 8526 8878 22159 8880
rect 5441 8875 5507 8878
rect 6821 8875 6887 8878
rect 0 8802 800 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 800 8742
rect 4061 8739 4127 8742
rect 4981 8802 5047 8805
rect 5390 8802 5396 8804
rect 4981 8800 5396 8802
rect 4981 8744 4986 8800
rect 5042 8744 5396 8800
rect 4981 8742 5396 8744
rect 4981 8739 5047 8742
rect 5390 8740 5396 8742
rect 5460 8740 5466 8804
rect 8342 8802 8402 8878
rect 22093 8875 22159 8878
rect 24853 8938 24919 8941
rect 26200 8938 27000 8968
rect 24853 8936 27000 8938
rect 24853 8880 24858 8936
rect 24914 8880 27000 8936
rect 24853 8878 27000 8880
rect 24853 8875 24919 8878
rect 26200 8848 27000 8878
rect 14406 8802 14412 8804
rect 8342 8742 14412 8802
rect 14406 8740 14412 8742
rect 14476 8740 14482 8804
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 5901 8666 5967 8669
rect 7230 8666 7236 8668
rect 5901 8664 7236 8666
rect 5901 8608 5906 8664
rect 5962 8608 7236 8664
rect 5901 8606 7236 8608
rect 5901 8603 5967 8606
rect 7230 8604 7236 8606
rect 7300 8604 7306 8668
rect 10225 8666 10291 8669
rect 12249 8666 12315 8669
rect 14038 8666 14044 8668
rect 10225 8664 12315 8666
rect 10225 8608 10230 8664
rect 10286 8608 12254 8664
rect 12310 8608 12315 8664
rect 10225 8606 12315 8608
rect 10225 8603 10291 8606
rect 12249 8603 12315 8606
rect 12390 8606 14044 8666
rect 2078 8530 2084 8532
rect 1996 8470 2084 8530
rect 2078 8468 2084 8470
rect 2148 8530 2154 8532
rect 5257 8530 5323 8533
rect 12390 8530 12450 8606
rect 14038 8604 14044 8606
rect 14108 8666 14114 8668
rect 15142 8666 15148 8668
rect 14108 8606 15148 8666
rect 14108 8604 14114 8606
rect 15142 8604 15148 8606
rect 15212 8604 15218 8668
rect 15694 8604 15700 8668
rect 15764 8666 15770 8668
rect 15764 8606 15946 8666
rect 15764 8604 15770 8606
rect 2148 8470 5090 8530
rect 2148 8468 2154 8470
rect 1945 8394 2011 8397
rect 2086 8394 2146 8468
rect 2681 8396 2747 8397
rect 2630 8394 2636 8396
rect 1945 8392 2146 8394
rect 1945 8336 1950 8392
rect 2006 8336 2146 8392
rect 1945 8334 2146 8336
rect 2590 8334 2636 8394
rect 2700 8392 2747 8396
rect 2742 8336 2747 8392
rect 1945 8331 2011 8334
rect 2630 8332 2636 8334
rect 2700 8332 2747 8336
rect 5030 8394 5090 8470
rect 5257 8528 12450 8530
rect 5257 8472 5262 8528
rect 5318 8472 12450 8528
rect 5257 8470 12450 8472
rect 5257 8467 5323 8470
rect 12750 8468 12756 8532
rect 12820 8530 12826 8532
rect 13261 8530 13327 8533
rect 12820 8528 13327 8530
rect 12820 8472 13266 8528
rect 13322 8472 13327 8528
rect 12820 8470 13327 8472
rect 12820 8468 12826 8470
rect 13261 8467 13327 8470
rect 14774 8468 14780 8532
rect 14844 8530 14850 8532
rect 15745 8530 15811 8533
rect 14844 8528 15811 8530
rect 14844 8472 15750 8528
rect 15806 8472 15811 8528
rect 14844 8470 15811 8472
rect 15886 8530 15946 8606
rect 20621 8530 20687 8533
rect 15886 8528 20687 8530
rect 15886 8472 20626 8528
rect 20682 8472 20687 8528
rect 15886 8470 20687 8472
rect 14844 8468 14850 8470
rect 15745 8467 15811 8470
rect 20621 8467 20687 8470
rect 15929 8394 15995 8397
rect 5030 8392 15995 8394
rect 5030 8336 15934 8392
rect 15990 8336 15995 8392
rect 5030 8334 15995 8336
rect 2681 8331 2747 8332
rect 15929 8331 15995 8334
rect 18505 8394 18571 8397
rect 18689 8394 18755 8397
rect 18505 8392 18755 8394
rect 18505 8336 18510 8392
rect 18566 8336 18694 8392
rect 18750 8336 18755 8392
rect 18505 8334 18755 8336
rect 18505 8331 18571 8334
rect 18689 8331 18755 8334
rect 4981 8258 5047 8261
rect 12014 8258 12020 8260
rect 4981 8256 12020 8258
rect 4981 8200 4986 8256
rect 5042 8200 12020 8256
rect 4981 8198 12020 8200
rect 4981 8195 5047 8198
rect 12014 8196 12020 8198
rect 12084 8196 12090 8260
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 3366 8060 3372 8124
rect 3436 8122 3442 8124
rect 3509 8122 3575 8125
rect 3436 8120 3575 8122
rect 3436 8064 3514 8120
rect 3570 8064 3575 8120
rect 3436 8062 3575 8064
rect 3436 8060 3442 8062
rect 3509 8059 3575 8062
rect 3969 8122 4035 8125
rect 7925 8122 7991 8125
rect 3969 8120 7991 8122
rect 3969 8064 3974 8120
rect 4030 8064 7930 8120
rect 7986 8064 7991 8120
rect 3969 8062 7991 8064
rect 3969 8059 4035 8062
rect 7925 8059 7991 8062
rect 8937 8122 9003 8125
rect 12801 8122 12867 8125
rect 8937 8120 12867 8122
rect 8937 8064 8942 8120
rect 8998 8064 12806 8120
rect 12862 8064 12867 8120
rect 8937 8062 12867 8064
rect 8937 8059 9003 8062
rect 12801 8059 12867 8062
rect 13537 8122 13603 8125
rect 13670 8122 13676 8124
rect 13537 8120 13676 8122
rect 13537 8064 13542 8120
rect 13598 8064 13676 8120
rect 13537 8062 13676 8064
rect 13537 8059 13603 8062
rect 13670 8060 13676 8062
rect 13740 8060 13746 8124
rect 13854 8060 13860 8124
rect 13924 8122 13930 8124
rect 14457 8122 14523 8125
rect 13924 8120 14523 8122
rect 13924 8064 14462 8120
rect 14518 8064 14523 8120
rect 13924 8062 14523 8064
rect 13924 8060 13930 8062
rect 14457 8059 14523 8062
rect 24853 8122 24919 8125
rect 26200 8122 27000 8152
rect 24853 8120 27000 8122
rect 24853 8064 24858 8120
rect 24914 8064 27000 8120
rect 24853 8062 27000 8064
rect 24853 8059 24919 8062
rect 26200 8032 27000 8062
rect 2405 7988 2471 7989
rect 1342 7924 1348 7988
rect 1412 7986 1418 7988
rect 2405 7986 2452 7988
rect 1412 7984 2452 7986
rect 1412 7928 2410 7984
rect 1412 7926 2452 7928
rect 1412 7924 1418 7926
rect 2405 7924 2452 7926
rect 2516 7924 2522 7988
rect 4429 7986 4495 7989
rect 17493 7986 17559 7989
rect 4429 7984 17559 7986
rect 4429 7928 4434 7984
rect 4490 7928 17498 7984
rect 17554 7928 17559 7984
rect 4429 7926 17559 7928
rect 2405 7923 2471 7924
rect 4429 7923 4495 7926
rect 17493 7923 17559 7926
rect 19609 7986 19675 7989
rect 20253 7986 20319 7989
rect 19609 7984 20319 7986
rect 19609 7928 19614 7984
rect 19670 7928 20258 7984
rect 20314 7928 20319 7984
rect 19609 7926 20319 7928
rect 19609 7923 19675 7926
rect 20253 7923 20319 7926
rect 7281 7850 7347 7853
rect 9581 7850 9647 7853
rect 20713 7850 20779 7853
rect 7281 7848 8402 7850
rect 7281 7792 7286 7848
rect 7342 7792 8402 7848
rect 7281 7790 8402 7792
rect 7281 7787 7347 7790
rect 1485 7714 1551 7717
rect 4889 7714 4955 7717
rect 1485 7712 4955 7714
rect 1485 7656 1490 7712
rect 1546 7656 4894 7712
rect 4950 7656 4955 7712
rect 1485 7654 4955 7656
rect 8342 7714 8402 7790
rect 9581 7848 20779 7850
rect 9581 7792 9586 7848
rect 9642 7792 20718 7848
rect 20774 7792 20779 7848
rect 9581 7790 20779 7792
rect 9581 7787 9647 7790
rect 20713 7787 20779 7790
rect 14273 7714 14339 7717
rect 8342 7712 14339 7714
rect 8342 7656 14278 7712
rect 14334 7656 14339 7712
rect 8342 7654 14339 7656
rect 1485 7651 1551 7654
rect 4889 7651 4955 7654
rect 14273 7651 14339 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 8569 7578 8635 7581
rect 8702 7578 8708 7580
rect 8569 7576 8708 7578
rect 8569 7520 8574 7576
rect 8630 7520 8708 7576
rect 8569 7518 8708 7520
rect 8569 7515 8635 7518
rect 8702 7516 8708 7518
rect 8772 7516 8778 7580
rect 11237 7578 11303 7581
rect 14222 7578 14228 7580
rect 11237 7576 14228 7578
rect 11237 7520 11242 7576
rect 11298 7520 14228 7576
rect 11237 7518 14228 7520
rect 11237 7515 11303 7518
rect 14222 7516 14228 7518
rect 14292 7516 14298 7580
rect 15142 7516 15148 7580
rect 15212 7578 15218 7580
rect 16481 7578 16547 7581
rect 15212 7576 16547 7578
rect 15212 7520 16486 7576
rect 16542 7520 16547 7576
rect 15212 7518 16547 7520
rect 15212 7516 15218 7518
rect 16481 7515 16547 7518
rect 4337 7444 4403 7445
rect 4286 7380 4292 7444
rect 4356 7442 4403 7444
rect 6821 7442 6887 7445
rect 22093 7442 22159 7445
rect 4356 7440 4448 7442
rect 4398 7384 4448 7440
rect 4356 7382 4448 7384
rect 6821 7440 22159 7442
rect 6821 7384 6826 7440
rect 6882 7384 22098 7440
rect 22154 7384 22159 7440
rect 6821 7382 22159 7384
rect 4356 7380 4403 7382
rect 4337 7379 4403 7380
rect 6821 7379 6887 7382
rect 22093 7379 22159 7382
rect 5901 7306 5967 7309
rect 23841 7306 23907 7309
rect 5901 7304 23907 7306
rect 5901 7248 5906 7304
rect 5962 7248 23846 7304
rect 23902 7248 23907 7304
rect 5901 7246 23907 7248
rect 5901 7243 5967 7246
rect 23841 7243 23907 7246
rect 24761 7306 24827 7309
rect 26200 7306 27000 7336
rect 24761 7304 27000 7306
rect 24761 7248 24766 7304
rect 24822 7248 27000 7304
rect 24761 7246 27000 7248
rect 24761 7243 24827 7246
rect 26200 7216 27000 7246
rect 4889 7170 4955 7173
rect 5022 7170 5028 7172
rect 4889 7168 5028 7170
rect 4889 7112 4894 7168
rect 4950 7112 5028 7168
rect 4889 7110 5028 7112
rect 4889 7107 4955 7110
rect 5022 7108 5028 7110
rect 5092 7108 5098 7172
rect 7005 7170 7071 7173
rect 7598 7170 7604 7172
rect 7005 7168 7604 7170
rect 7005 7112 7010 7168
rect 7066 7112 7604 7168
rect 7005 7110 7604 7112
rect 7005 7107 7071 7110
rect 7598 7108 7604 7110
rect 7668 7108 7674 7172
rect 13486 7108 13492 7172
rect 13556 7170 13562 7172
rect 19333 7170 19399 7173
rect 19885 7170 19951 7173
rect 13556 7168 19951 7170
rect 13556 7112 19338 7168
rect 19394 7112 19890 7168
rect 19946 7112 19951 7168
rect 13556 7110 19951 7112
rect 13556 7108 13562 7110
rect 19333 7107 19399 7110
rect 19885 7107 19951 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 4889 7034 4955 7037
rect 6453 7034 6519 7037
rect 4889 7032 6519 7034
rect 4889 6976 4894 7032
rect 4950 6976 6458 7032
rect 6514 6976 6519 7032
rect 4889 6974 6519 6976
rect 4889 6971 4955 6974
rect 6453 6971 6519 6974
rect 6637 7034 6703 7037
rect 17585 7034 17651 7037
rect 6637 7032 12818 7034
rect 6637 6976 6642 7032
rect 6698 6976 12818 7032
rect 6637 6974 12818 6976
rect 6637 6971 6703 6974
rect 7097 6898 7163 6901
rect 8569 6898 8635 6901
rect 7097 6896 8635 6898
rect 7097 6840 7102 6896
rect 7158 6840 8574 6896
rect 8630 6840 8635 6896
rect 7097 6838 8635 6840
rect 7097 6835 7163 6838
rect 8569 6835 8635 6838
rect 11329 6898 11395 6901
rect 12341 6898 12407 6901
rect 12617 6900 12683 6901
rect 12566 6898 12572 6900
rect 11329 6896 12407 6898
rect 11329 6840 11334 6896
rect 11390 6840 12346 6896
rect 12402 6840 12407 6896
rect 11329 6838 12407 6840
rect 12526 6838 12572 6898
rect 12636 6896 12683 6900
rect 12678 6840 12683 6896
rect 11329 6835 11395 6838
rect 12341 6835 12407 6838
rect 12566 6836 12572 6838
rect 12636 6836 12683 6840
rect 12758 6898 12818 6974
rect 13494 7032 17651 7034
rect 13494 6976 17590 7032
rect 17646 6976 17651 7032
rect 13494 6974 17651 6976
rect 13494 6898 13554 6974
rect 17585 6971 17651 6974
rect 12758 6838 13554 6898
rect 14917 6898 14983 6901
rect 15929 6898 15995 6901
rect 14917 6896 15995 6898
rect 14917 6840 14922 6896
rect 14978 6840 15934 6896
rect 15990 6840 15995 6896
rect 14917 6838 15995 6840
rect 12617 6835 12683 6836
rect 14917 6835 14983 6838
rect 15929 6835 15995 6838
rect 16481 6898 16547 6901
rect 17585 6898 17651 6901
rect 16481 6896 17651 6898
rect 16481 6840 16486 6896
rect 16542 6840 17590 6896
rect 17646 6840 17651 6896
rect 16481 6838 17651 6840
rect 16481 6835 16547 6838
rect 17585 6835 17651 6838
rect 18229 6898 18295 6901
rect 24669 6898 24735 6901
rect 18229 6896 24735 6898
rect 18229 6840 18234 6896
rect 18290 6840 24674 6896
rect 24730 6840 24735 6896
rect 18229 6838 24735 6840
rect 18229 6835 18295 6838
rect 24669 6835 24735 6838
rect 4061 6762 4127 6765
rect 2730 6760 4127 6762
rect 2730 6704 4066 6760
rect 4122 6704 4127 6760
rect 2730 6702 4127 6704
rect 0 6490 800 6520
rect 2730 6490 2790 6702
rect 4061 6699 4127 6702
rect 5390 6700 5396 6764
rect 5460 6762 5466 6764
rect 20069 6762 20135 6765
rect 5460 6760 20135 6762
rect 5460 6704 20074 6760
rect 20130 6704 20135 6760
rect 5460 6702 20135 6704
rect 5460 6700 5466 6702
rect 20069 6699 20135 6702
rect 8569 6626 8635 6629
rect 14733 6626 14799 6629
rect 8569 6624 14799 6626
rect 8569 6568 8574 6624
rect 8630 6568 14738 6624
rect 14794 6568 14799 6624
rect 8569 6566 14799 6568
rect 8569 6563 8635 6566
rect 14733 6563 14799 6566
rect 14917 6626 14983 6629
rect 15469 6626 15535 6629
rect 15837 6626 15903 6629
rect 14917 6624 15903 6626
rect 14917 6568 14922 6624
rect 14978 6568 15474 6624
rect 15530 6568 15842 6624
rect 15898 6568 15903 6624
rect 14917 6566 15903 6568
rect 14917 6563 14983 6566
rect 15469 6563 15535 6566
rect 15837 6563 15903 6566
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 0 6430 2790 6490
rect 0 6400 800 6430
rect 11094 6428 11100 6492
rect 11164 6490 11170 6492
rect 12525 6490 12591 6493
rect 13537 6492 13603 6493
rect 13486 6490 13492 6492
rect 11164 6488 12591 6490
rect 11164 6432 12530 6488
rect 12586 6432 12591 6488
rect 11164 6430 12591 6432
rect 13446 6430 13492 6490
rect 13556 6488 13603 6492
rect 15469 6492 15535 6493
rect 15469 6490 15516 6492
rect 13598 6432 13603 6488
rect 11164 6428 11170 6430
rect 12525 6427 12591 6430
rect 13486 6428 13492 6430
rect 13556 6428 13603 6432
rect 15424 6488 15516 6490
rect 15424 6432 15474 6488
rect 15424 6430 15516 6432
rect 13537 6427 13603 6428
rect 15469 6428 15516 6430
rect 15580 6428 15586 6492
rect 15837 6490 15903 6493
rect 16757 6490 16823 6493
rect 15837 6488 16823 6490
rect 15837 6432 15842 6488
rect 15898 6432 16762 6488
rect 16818 6432 16823 6488
rect 15837 6430 16823 6432
rect 15469 6427 15535 6428
rect 15837 6427 15903 6430
rect 16757 6427 16823 6430
rect 25037 6490 25103 6493
rect 26200 6490 27000 6520
rect 25037 6488 27000 6490
rect 25037 6432 25042 6488
rect 25098 6432 27000 6488
rect 25037 6430 27000 6432
rect 25037 6427 25103 6430
rect 26200 6400 27000 6430
rect 5073 6354 5139 6357
rect 22093 6354 22159 6357
rect 5073 6352 22159 6354
rect 5073 6296 5078 6352
rect 5134 6296 22098 6352
rect 22154 6296 22159 6352
rect 5073 6294 22159 6296
rect 5073 6291 5139 6294
rect 22093 6291 22159 6294
rect 4337 6218 4403 6221
rect 20805 6218 20871 6221
rect 4337 6216 20871 6218
rect 4337 6160 4342 6216
rect 4398 6160 20810 6216
rect 20866 6160 20871 6216
rect 4337 6158 20871 6160
rect 4337 6155 4403 6158
rect 20805 6155 20871 6158
rect 12157 6082 12223 6085
rect 12617 6082 12683 6085
rect 12157 6080 12683 6082
rect 12157 6024 12162 6080
rect 12218 6024 12622 6080
rect 12678 6024 12683 6080
rect 12157 6022 12683 6024
rect 12157 6019 12223 6022
rect 12617 6019 12683 6022
rect 14958 6020 14964 6084
rect 15028 6082 15034 6084
rect 16757 6082 16823 6085
rect 19609 6082 19675 6085
rect 15028 6080 19675 6082
rect 15028 6024 16762 6080
rect 16818 6024 19614 6080
rect 19670 6024 19675 6080
rect 15028 6022 19675 6024
rect 15028 6020 15034 6022
rect 16757 6019 16823 6022
rect 19609 6019 19675 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 5165 5946 5231 5949
rect 11830 5946 11836 5948
rect 5165 5944 11836 5946
rect 5165 5888 5170 5944
rect 5226 5888 11836 5944
rect 5165 5886 11836 5888
rect 5165 5883 5231 5886
rect 11830 5884 11836 5886
rect 11900 5884 11906 5948
rect 11973 5946 12039 5949
rect 12341 5946 12407 5949
rect 11973 5944 12407 5946
rect 11973 5888 11978 5944
rect 12034 5888 12346 5944
rect 12402 5888 12407 5944
rect 11973 5886 12407 5888
rect 11973 5883 12039 5886
rect 12341 5883 12407 5886
rect 13537 5946 13603 5949
rect 17125 5946 17191 5949
rect 13537 5944 17191 5946
rect 13537 5888 13542 5944
rect 13598 5888 17130 5944
rect 17186 5888 17191 5944
rect 13537 5886 17191 5888
rect 13537 5883 13603 5886
rect 17125 5883 17191 5886
rect 18137 5946 18203 5949
rect 19333 5946 19399 5949
rect 19701 5946 19767 5949
rect 18137 5944 19767 5946
rect 18137 5888 18142 5944
rect 18198 5888 19338 5944
rect 19394 5888 19706 5944
rect 19762 5888 19767 5944
rect 18137 5886 19767 5888
rect 18137 5883 18203 5886
rect 19333 5883 19399 5886
rect 19701 5883 19767 5886
rect 7649 5810 7715 5813
rect 14774 5810 14780 5812
rect 7649 5808 14780 5810
rect 7649 5752 7654 5808
rect 7710 5752 14780 5808
rect 7649 5750 14780 5752
rect 7649 5747 7715 5750
rect 14774 5748 14780 5750
rect 14844 5748 14850 5812
rect 15142 5748 15148 5812
rect 15212 5810 15218 5812
rect 15561 5810 15627 5813
rect 15212 5808 15627 5810
rect 15212 5752 15566 5808
rect 15622 5752 15627 5808
rect 15212 5750 15627 5752
rect 15212 5748 15218 5750
rect 15561 5747 15627 5750
rect 4153 5676 4219 5677
rect 4102 5674 4108 5676
rect 4062 5614 4108 5674
rect 4172 5672 4219 5676
rect 4214 5616 4219 5672
rect 4102 5612 4108 5614
rect 4172 5612 4219 5616
rect 4153 5611 4219 5612
rect 7281 5674 7347 5677
rect 7925 5674 7991 5677
rect 7281 5672 7991 5674
rect 7281 5616 7286 5672
rect 7342 5616 7930 5672
rect 7986 5616 7991 5672
rect 7281 5614 7991 5616
rect 7281 5611 7347 5614
rect 7925 5611 7991 5614
rect 8753 5674 8819 5677
rect 9070 5674 9076 5676
rect 8753 5672 9076 5674
rect 8753 5616 8758 5672
rect 8814 5616 9076 5672
rect 8753 5614 9076 5616
rect 8753 5611 8819 5614
rect 9070 5612 9076 5614
rect 9140 5674 9146 5676
rect 24577 5674 24643 5677
rect 9140 5672 24643 5674
rect 9140 5616 24582 5672
rect 24638 5616 24643 5672
rect 9140 5614 24643 5616
rect 9140 5612 9146 5614
rect 24577 5611 24643 5614
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 1301 5538 1367 5541
rect 7557 5538 7623 5541
rect 1301 5536 7623 5538
rect 1301 5480 1306 5536
rect 1362 5480 7562 5536
rect 7618 5480 7623 5536
rect 1301 5478 7623 5480
rect 1301 5475 1367 5478
rect 7557 5475 7623 5478
rect 11881 5538 11947 5541
rect 14733 5538 14799 5541
rect 11881 5536 14799 5538
rect 11881 5480 11886 5536
rect 11942 5480 14738 5536
rect 14794 5480 14799 5536
rect 11881 5478 14799 5480
rect 11881 5475 11947 5478
rect 14733 5475 14799 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 5717 5402 5783 5405
rect 7649 5402 7715 5405
rect 14917 5402 14983 5405
rect 16665 5402 16731 5405
rect 5717 5400 7715 5402
rect 5717 5344 5722 5400
rect 5778 5344 7654 5400
rect 7710 5344 7715 5400
rect 5717 5342 7715 5344
rect 5717 5339 5783 5342
rect 7649 5339 7715 5342
rect 10964 5400 16731 5402
rect 10964 5344 14922 5400
rect 14978 5344 16670 5400
rect 16726 5344 16731 5400
rect 10964 5342 16731 5344
rect 10964 5269 11024 5342
rect 14917 5339 14983 5342
rect 16665 5339 16731 5342
rect 7649 5266 7715 5269
rect 10961 5266 11027 5269
rect 7649 5264 11027 5266
rect 7649 5208 7654 5264
rect 7710 5208 10966 5264
rect 11022 5208 11027 5264
rect 7649 5206 11027 5208
rect 7649 5203 7715 5206
rect 10961 5203 11027 5206
rect 12014 5204 12020 5268
rect 12084 5266 12090 5268
rect 23933 5266 23999 5269
rect 12084 5264 23999 5266
rect 12084 5208 23938 5264
rect 23994 5208 23999 5264
rect 12084 5206 23999 5208
rect 12084 5204 12090 5206
rect 23933 5203 23999 5206
rect 9305 5130 9371 5133
rect 18413 5130 18479 5133
rect 19977 5130 20043 5133
rect 9305 5128 20043 5130
rect 9305 5072 9310 5128
rect 9366 5072 18418 5128
rect 18474 5072 19982 5128
rect 20038 5072 20043 5128
rect 9305 5070 20043 5072
rect 9305 5067 9371 5070
rect 18413 5067 18479 5070
rect 19977 5067 20043 5070
rect 3918 4932 3924 4996
rect 3988 4994 3994 4996
rect 9121 4994 9187 4997
rect 3988 4992 9187 4994
rect 3988 4936 9126 4992
rect 9182 4936 9187 4992
rect 3988 4934 9187 4936
rect 3988 4932 3994 4934
rect 9121 4931 9187 4934
rect 13905 4994 13971 4997
rect 19241 4994 19307 4997
rect 13905 4992 19307 4994
rect 13905 4936 13910 4992
rect 13966 4936 19246 4992
rect 19302 4936 19307 4992
rect 13905 4934 19307 4936
rect 13905 4931 13971 4934
rect 19241 4931 19307 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 5625 4858 5691 4861
rect 9806 4858 9812 4860
rect 5625 4856 9812 4858
rect 5625 4800 5630 4856
rect 5686 4800 9812 4856
rect 5625 4798 9812 4800
rect 5625 4795 5691 4798
rect 9806 4796 9812 4798
rect 9876 4858 9882 4860
rect 12341 4858 12407 4861
rect 9876 4856 12407 4858
rect 9876 4800 12346 4856
rect 12402 4800 12407 4856
rect 9876 4798 12407 4800
rect 9876 4796 9882 4798
rect 12341 4795 12407 4798
rect 14273 4858 14339 4861
rect 21173 4860 21239 4861
rect 21173 4858 21220 4860
rect 14273 4856 21220 4858
rect 21284 4858 21290 4860
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 14273 4800 14278 4856
rect 14334 4800 21178 4856
rect 14273 4798 21220 4800
rect 14273 4795 14339 4798
rect 21173 4796 21220 4798
rect 21284 4798 21366 4858
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 21284 4796 21290 4798
rect 21173 4795 21239 4796
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 3233 4722 3299 4725
rect 8293 4722 8359 4725
rect 3233 4720 8359 4722
rect 3233 4664 3238 4720
rect 3294 4664 8298 4720
rect 8354 4664 8359 4720
rect 3233 4662 8359 4664
rect 3233 4659 3299 4662
rect 8293 4659 8359 4662
rect 11830 4660 11836 4724
rect 11900 4722 11906 4724
rect 20713 4722 20779 4725
rect 11900 4720 20779 4722
rect 11900 4664 20718 4720
rect 20774 4664 20779 4720
rect 11900 4662 20779 4664
rect 11900 4660 11906 4662
rect 20713 4659 20779 4662
rect 1669 4586 1735 4589
rect 11789 4586 11855 4589
rect 1669 4584 11855 4586
rect 1669 4528 1674 4584
rect 1730 4528 11794 4584
rect 11850 4528 11855 4584
rect 1669 4526 11855 4528
rect 1669 4523 1735 4526
rect 11789 4523 11855 4526
rect 12341 4586 12407 4589
rect 22645 4586 22711 4589
rect 12341 4584 22711 4586
rect 12341 4528 12346 4584
rect 12402 4528 22650 4584
rect 22706 4528 22711 4584
rect 12341 4526 22711 4528
rect 12341 4523 12407 4526
rect 22645 4523 22711 4526
rect 8477 4452 8543 4453
rect 8477 4448 8524 4452
rect 8588 4450 8594 4452
rect 13854 4450 13860 4452
rect 8477 4392 8482 4448
rect 8477 4388 8524 4392
rect 8588 4390 8634 4450
rect 8710 4390 13860 4450
rect 8588 4388 8594 4390
rect 8477 4387 8543 4388
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 4061 4314 4127 4317
rect 2730 4312 4127 4314
rect 2730 4256 4066 4312
rect 4122 4256 4127 4312
rect 2730 4254 4127 4256
rect 0 4178 800 4208
rect 2730 4178 2790 4254
rect 4061 4251 4127 4254
rect 8385 4314 8451 4317
rect 8710 4314 8770 4390
rect 13854 4388 13860 4390
rect 13924 4388 13930 4452
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 8385 4312 8770 4314
rect 8385 4256 8390 4312
rect 8446 4256 8770 4312
rect 8385 4254 8770 4256
rect 8845 4314 8911 4317
rect 8845 4312 15210 4314
rect 8845 4256 8850 4312
rect 8906 4256 15210 4312
rect 8845 4254 15210 4256
rect 8385 4251 8451 4254
rect 8845 4251 8911 4254
rect 0 4118 2790 4178
rect 2865 4178 2931 4181
rect 9673 4178 9739 4181
rect 2865 4176 9739 4178
rect 2865 4120 2870 4176
rect 2926 4120 9678 4176
rect 9734 4120 9739 4176
rect 2865 4118 9739 4120
rect 0 4088 800 4118
rect 2865 4115 2931 4118
rect 9673 4115 9739 4118
rect 1669 4044 1735 4045
rect 1669 4040 1716 4044
rect 1780 4042 1786 4044
rect 2865 4042 2931 4045
rect 3550 4042 3556 4044
rect 1669 3984 1674 4040
rect 1669 3980 1716 3984
rect 1780 3982 1826 4042
rect 2865 4040 3556 4042
rect 2865 3984 2870 4040
rect 2926 3984 3556 4040
rect 2865 3982 3556 3984
rect 1780 3980 1786 3982
rect 1669 3979 1735 3980
rect 2865 3979 2931 3982
rect 3550 3980 3556 3982
rect 3620 3980 3626 4044
rect 5574 3980 5580 4044
rect 5644 4042 5650 4044
rect 5901 4042 5967 4045
rect 5644 4040 5967 4042
rect 5644 3984 5906 4040
rect 5962 3984 5967 4040
rect 5644 3982 5967 3984
rect 5644 3980 5650 3982
rect 5901 3979 5967 3982
rect 6085 4042 6151 4045
rect 12617 4042 12683 4045
rect 6085 4040 12683 4042
rect 6085 3984 6090 4040
rect 6146 3984 12622 4040
rect 12678 3984 12683 4040
rect 6085 3982 12683 3984
rect 15150 4042 15210 4254
rect 17166 4116 17172 4180
rect 17236 4178 17242 4180
rect 19425 4178 19491 4181
rect 17236 4176 19491 4178
rect 17236 4120 19430 4176
rect 19486 4120 19491 4176
rect 17236 4118 19491 4120
rect 17236 4116 17242 4118
rect 19425 4115 19491 4118
rect 18045 4042 18111 4045
rect 15150 4040 18111 4042
rect 15150 3984 18050 4040
rect 18106 3984 18111 4040
rect 15150 3982 18111 3984
rect 6085 3979 6151 3982
rect 12617 3979 12683 3982
rect 18045 3979 18111 3982
rect 19006 3980 19012 4044
rect 19076 4042 19082 4044
rect 19701 4042 19767 4045
rect 19076 4040 19767 4042
rect 19076 3984 19706 4040
rect 19762 3984 19767 4040
rect 19076 3982 19767 3984
rect 19076 3980 19082 3982
rect 19701 3979 19767 3982
rect 20478 3980 20484 4044
rect 20548 4042 20554 4044
rect 20621 4042 20687 4045
rect 20548 4040 20687 4042
rect 20548 3984 20626 4040
rect 20682 3984 20687 4040
rect 20548 3982 20687 3984
rect 20548 3980 20554 3982
rect 20621 3979 20687 3982
rect 23381 4042 23447 4045
rect 26200 4042 27000 4072
rect 23381 4040 27000 4042
rect 23381 3984 23386 4040
rect 23442 3984 27000 4040
rect 23381 3982 27000 3984
rect 23381 3979 23447 3982
rect 26200 3952 27000 3982
rect 13445 3906 13511 3909
rect 19885 3906 19951 3909
rect 13445 3904 19951 3906
rect 13445 3848 13450 3904
rect 13506 3848 19890 3904
rect 19946 3848 19951 3904
rect 13445 3846 19951 3848
rect 13445 3843 13511 3846
rect 19885 3843 19951 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 4613 3770 4679 3773
rect 11053 3770 11119 3773
rect 4613 3768 11119 3770
rect 4613 3712 4618 3768
rect 4674 3712 11058 3768
rect 11114 3712 11119 3768
rect 4613 3710 11119 3712
rect 4613 3707 4679 3710
rect 11053 3707 11119 3710
rect 14457 3770 14523 3773
rect 15326 3770 15332 3772
rect 14457 3768 15332 3770
rect 14457 3712 14462 3768
rect 14518 3712 15332 3768
rect 14457 3710 15332 3712
rect 14457 3707 14523 3710
rect 15326 3708 15332 3710
rect 15396 3708 15402 3772
rect 24209 3770 24275 3773
rect 24526 3770 24532 3772
rect 24209 3768 24532 3770
rect 24209 3712 24214 3768
rect 24270 3712 24532 3768
rect 24209 3710 24532 3712
rect 24209 3707 24275 3710
rect 24526 3708 24532 3710
rect 24596 3708 24602 3772
rect 6637 3634 6703 3637
rect 7782 3634 7788 3636
rect 6637 3632 7788 3634
rect 6637 3576 6642 3632
rect 6698 3576 7788 3632
rect 6637 3574 7788 3576
rect 6637 3571 6703 3574
rect 7782 3572 7788 3574
rect 7852 3572 7858 3636
rect 7925 3634 7991 3637
rect 17769 3634 17835 3637
rect 7925 3632 17835 3634
rect 7925 3576 7930 3632
rect 7986 3576 17774 3632
rect 17830 3576 17835 3632
rect 7925 3574 17835 3576
rect 7925 3571 7991 3574
rect 17769 3571 17835 3574
rect 22318 3572 22324 3636
rect 22388 3634 22394 3636
rect 23841 3634 23907 3637
rect 22388 3632 23907 3634
rect 22388 3576 23846 3632
rect 23902 3576 23907 3632
rect 22388 3574 23907 3576
rect 22388 3572 22394 3574
rect 23841 3571 23907 3574
rect 7465 3498 7531 3501
rect 14958 3498 14964 3500
rect 7465 3496 14964 3498
rect 7465 3440 7470 3496
rect 7526 3440 14964 3496
rect 7465 3438 14964 3440
rect 7465 3435 7531 3438
rect 14958 3436 14964 3438
rect 15028 3436 15034 3500
rect 2681 3362 2747 3365
rect 7649 3362 7715 3365
rect 2681 3360 7715 3362
rect 2681 3304 2686 3360
rect 2742 3304 7654 3360
rect 7710 3304 7715 3360
rect 2681 3302 7715 3304
rect 2681 3299 2747 3302
rect 7649 3299 7715 3302
rect 8753 3362 8819 3365
rect 10910 3362 10916 3364
rect 8753 3360 10916 3362
rect 8753 3304 8758 3360
rect 8814 3304 10916 3360
rect 8753 3302 10916 3304
rect 8753 3299 8819 3302
rect 10910 3300 10916 3302
rect 10980 3362 10986 3364
rect 15101 3362 15167 3365
rect 10980 3360 15167 3362
rect 10980 3304 15106 3360
rect 15162 3304 15167 3360
rect 10980 3302 15167 3304
rect 10980 3300 10986 3302
rect 15101 3299 15167 3302
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 1853 3226 1919 3229
rect 7649 3226 7715 3229
rect 14590 3226 14596 3228
rect 1853 3224 7715 3226
rect 1853 3168 1858 3224
rect 1914 3168 7654 3224
rect 7710 3168 7715 3224
rect 1853 3166 7715 3168
rect 1853 3163 1919 3166
rect 7649 3163 7715 3166
rect 12390 3166 14596 3226
rect 3877 3090 3943 3093
rect 12390 3090 12450 3166
rect 14590 3164 14596 3166
rect 14660 3164 14666 3228
rect 22277 3226 22343 3229
rect 26200 3226 27000 3256
rect 22277 3224 27000 3226
rect 22277 3168 22282 3224
rect 22338 3168 27000 3224
rect 22277 3166 27000 3168
rect 22277 3163 22343 3166
rect 26200 3136 27000 3166
rect 3877 3088 12450 3090
rect 3877 3032 3882 3088
rect 3938 3032 12450 3088
rect 3877 3030 12450 3032
rect 3877 3027 3943 3030
rect 14406 3028 14412 3092
rect 14476 3090 14482 3092
rect 22093 3090 22159 3093
rect 14476 3088 22159 3090
rect 14476 3032 22098 3088
rect 22154 3032 22159 3088
rect 14476 3030 22159 3032
rect 14476 3028 14482 3030
rect 22093 3027 22159 3030
rect 6177 2954 6243 2957
rect 6494 2954 6500 2956
rect 6177 2952 6500 2954
rect 6177 2896 6182 2952
rect 6238 2896 6500 2952
rect 6177 2894 6500 2896
rect 6177 2891 6243 2894
rect 6494 2892 6500 2894
rect 6564 2892 6570 2956
rect 8937 2954 9003 2957
rect 18505 2954 18571 2957
rect 8937 2952 18571 2954
rect 8937 2896 8942 2952
rect 8998 2896 18510 2952
rect 18566 2896 18571 2952
rect 8937 2894 18571 2896
rect 8937 2891 9003 2894
rect 18505 2891 18571 2894
rect 18873 2954 18939 2957
rect 19149 2954 19215 2957
rect 18873 2952 19215 2954
rect 18873 2896 18878 2952
rect 18934 2896 19154 2952
rect 19210 2896 19215 2952
rect 18873 2894 19215 2896
rect 18873 2891 18939 2894
rect 19149 2891 19215 2894
rect 8293 2818 8359 2821
rect 9254 2818 9260 2820
rect 8293 2816 9260 2818
rect 8293 2760 8298 2816
rect 8354 2760 9260 2816
rect 8293 2758 9260 2760
rect 8293 2755 8359 2758
rect 9254 2756 9260 2758
rect 9324 2756 9330 2820
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 7230 2620 7236 2684
rect 7300 2682 7306 2684
rect 8385 2682 8451 2685
rect 7300 2680 8451 2682
rect 7300 2624 8390 2680
rect 8446 2624 8451 2680
rect 7300 2622 8451 2624
rect 7300 2620 7306 2622
rect 8385 2619 8451 2622
rect 5441 2546 5507 2549
rect 14089 2546 14155 2549
rect 5441 2544 14155 2546
rect 5441 2488 5446 2544
rect 5502 2488 14094 2544
rect 14150 2488 14155 2544
rect 5441 2486 14155 2488
rect 5441 2483 5507 2486
rect 14089 2483 14155 2486
rect 6361 2410 6427 2413
rect 17861 2410 17927 2413
rect 6361 2408 17927 2410
rect 6361 2352 6366 2408
rect 6422 2352 17866 2408
rect 17922 2352 17927 2408
rect 6361 2350 17927 2352
rect 6361 2347 6427 2350
rect 17861 2347 17927 2350
rect 22185 2410 22251 2413
rect 26200 2410 27000 2440
rect 22185 2408 27000 2410
rect 22185 2352 22190 2408
rect 22246 2352 27000 2408
rect 22185 2350 27000 2352
rect 22185 2347 22251 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 8385 2138 8451 2141
rect 8385 2136 16590 2138
rect 8385 2080 8390 2136
rect 8446 2080 16590 2136
rect 8385 2078 16590 2080
rect 8385 2075 8451 2078
rect 13537 2002 13603 2005
rect 6870 2000 13603 2002
rect 6870 1944 13542 2000
rect 13598 1944 13603 2000
rect 6870 1942 13603 1944
rect 16530 2002 16590 2078
rect 20345 2002 20411 2005
rect 16530 2000 20411 2002
rect 16530 1944 20350 2000
rect 20406 1944 20411 2000
rect 16530 1942 20411 1944
rect 0 1866 800 1896
rect 4654 1866 4660 1868
rect 0 1806 4660 1866
rect 0 1776 800 1806
rect 4654 1804 4660 1806
rect 4724 1804 4730 1868
rect 2313 1730 2379 1733
rect 6870 1730 6930 1942
rect 13537 1939 13603 1942
rect 20345 1939 20411 1942
rect 8886 1804 8892 1868
rect 8956 1866 8962 1868
rect 21633 1866 21699 1869
rect 8956 1864 21699 1866
rect 8956 1808 21638 1864
rect 21694 1808 21699 1864
rect 8956 1806 21699 1808
rect 8956 1804 8962 1806
rect 21633 1803 21699 1806
rect 2313 1728 6930 1730
rect 2313 1672 2318 1728
rect 2374 1672 6930 1728
rect 2313 1670 6930 1672
rect 12525 1730 12591 1733
rect 20846 1730 20852 1732
rect 12525 1728 20852 1730
rect 12525 1672 12530 1728
rect 12586 1672 20852 1728
rect 12525 1670 20852 1672
rect 2313 1667 2379 1670
rect 12525 1667 12591 1670
rect 20846 1668 20852 1670
rect 20916 1668 20922 1732
rect 4470 1532 4476 1596
rect 4540 1594 4546 1596
rect 15142 1594 15148 1596
rect 4540 1534 15148 1594
rect 4540 1532 4546 1534
rect 15142 1532 15148 1534
rect 15212 1532 15218 1596
rect 22277 1594 22343 1597
rect 26200 1594 27000 1624
rect 22277 1592 27000 1594
rect 22277 1536 22282 1592
rect 22338 1536 27000 1592
rect 22277 1534 27000 1536
rect 22277 1531 22343 1534
rect 26200 1504 27000 1534
rect 6821 1458 6887 1461
rect 15285 1458 15351 1461
rect 6821 1456 15351 1458
rect 6821 1400 6826 1456
rect 6882 1400 15290 1456
rect 15346 1400 15351 1456
rect 6821 1398 15351 1400
rect 6821 1395 6887 1398
rect 15285 1395 15351 1398
rect 7598 1260 7604 1324
rect 7668 1322 7674 1324
rect 7925 1322 7991 1325
rect 7668 1320 7991 1322
rect 7668 1264 7930 1320
rect 7986 1264 7991 1320
rect 7668 1262 7991 1264
rect 7668 1260 7674 1262
rect 7925 1259 7991 1262
rect 17033 1322 17099 1325
rect 19006 1322 19012 1324
rect 17033 1320 19012 1322
rect 17033 1264 17038 1320
rect 17094 1264 19012 1320
rect 17033 1262 19012 1264
rect 17033 1259 17099 1262
rect 19006 1260 19012 1262
rect 19076 1260 19082 1324
rect 5022 1124 5028 1188
rect 5092 1186 5098 1188
rect 17401 1186 17467 1189
rect 5092 1184 17467 1186
rect 5092 1128 17406 1184
rect 17462 1128 17467 1184
rect 5092 1126 17467 1128
rect 5092 1124 5098 1126
rect 17401 1123 17467 1126
rect 17534 1124 17540 1188
rect 17604 1186 17610 1188
rect 23289 1186 23355 1189
rect 17604 1184 23355 1186
rect 17604 1128 23294 1184
rect 23350 1128 23355 1184
rect 17604 1126 23355 1128
rect 17604 1124 17610 1126
rect 23289 1123 23355 1126
rect 7782 988 7788 1052
rect 7852 1050 7858 1052
rect 16982 1050 16988 1052
rect 7852 990 16988 1050
rect 7852 988 7858 990
rect 16982 988 16988 990
rect 17052 988 17058 1052
rect 20805 1050 20871 1053
rect 17174 1048 20871 1050
rect 17174 992 20810 1048
rect 20866 992 20871 1048
rect 17174 990 20871 992
rect 2630 852 2636 916
rect 2700 914 2706 916
rect 17033 914 17099 917
rect 2700 912 17099 914
rect 2700 856 17038 912
rect 17094 856 17099 912
rect 2700 854 17099 856
rect 2700 852 2706 854
rect 17033 851 17099 854
rect 1342 716 1348 780
rect 1412 778 1418 780
rect 17174 778 17234 990
rect 20805 987 20871 990
rect 18689 914 18755 917
rect 1412 718 17234 778
rect 17358 912 18755 914
rect 17358 856 18694 912
rect 18750 856 18755 912
rect 17358 854 18755 856
rect 1412 716 1418 718
rect 1158 580 1164 644
rect 1228 642 1234 644
rect 17358 642 17418 854
rect 18689 851 18755 854
rect 24945 778 25011 781
rect 26200 778 27000 808
rect 24945 776 27000 778
rect 24945 720 24950 776
rect 25006 720 27000 776
rect 24945 718 27000 720
rect 24945 715 25011 718
rect 26200 688 27000 718
rect 1228 582 17418 642
rect 1228 580 1234 582
rect 974 444 980 508
rect 1044 506 1050 508
rect 16297 506 16363 509
rect 1044 504 16363 506
rect 1044 448 16302 504
rect 16358 448 16363 504
rect 1044 446 16363 448
rect 1044 444 1050 446
rect 16297 443 16363 446
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 21036 47636 21100 47700
rect 16252 47500 16316 47564
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 20484 46956 20548 47020
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 15332 42604 15396 42668
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 12204 41516 12268 41580
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 19748 40020 19812 40084
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 16436 35804 16500 35868
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 15700 34444 15764 34508
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 18644 30832 18708 30836
rect 18644 30776 18658 30832
rect 18658 30776 18708 30832
rect 18644 30772 18708 30776
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 22692 29004 22756 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 18644 27508 18708 27572
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 17724 26420 17788 26484
rect 19012 26344 19076 26348
rect 19012 26288 19026 26344
rect 19026 26288 19076 26344
rect 19012 26284 19076 26288
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 11652 25740 11716 25804
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 16252 25332 16316 25396
rect 21036 25332 21100 25396
rect 24716 25332 24780 25396
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 20852 24984 20916 24988
rect 20852 24928 20866 24984
rect 20866 24928 20916 24984
rect 20852 24924 20916 24928
rect 22140 24924 22204 24988
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 13492 23428 13556 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 24532 22612 24596 22676
rect 10916 22476 10980 22540
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 4660 21524 4724 21588
rect 20484 21388 20548 21452
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 17540 21116 17604 21180
rect 12572 20844 12636 20908
rect 14228 20768 14292 20772
rect 14228 20712 14242 20768
rect 14242 20712 14292 20768
rect 14228 20708 14292 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 14964 19620 15028 19684
rect 20668 19680 20732 19684
rect 20668 19624 20682 19680
rect 20682 19624 20732 19680
rect 20668 19620 20732 19624
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 15148 19348 15212 19412
rect 16988 19076 17052 19140
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 14964 18940 15028 19004
rect 21036 18940 21100 19004
rect 15148 18804 15212 18868
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 3556 18260 3620 18324
rect 9260 18048 9324 18052
rect 9260 17992 9274 18048
rect 9274 17992 9324 18048
rect 9260 17988 9324 17992
rect 11836 18048 11900 18052
rect 11836 17992 11850 18048
rect 11850 17992 11900 18048
rect 11836 17988 11900 17992
rect 12020 18048 12084 18052
rect 12020 17992 12034 18048
rect 12034 17992 12084 18048
rect 12020 17988 12084 17992
rect 14044 17988 14108 18052
rect 15884 17988 15948 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 15700 17912 15764 17916
rect 15700 17856 15750 17912
rect 15750 17856 15764 17912
rect 15700 17852 15764 17856
rect 22324 17852 22388 17916
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 22692 17308 22756 17372
rect 4292 16900 4356 16964
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 6500 16688 6564 16692
rect 6500 16632 6514 16688
rect 6514 16632 6564 16688
rect 6500 16628 6564 16632
rect 8340 16688 8404 16692
rect 8340 16632 8354 16688
rect 8354 16632 8404 16688
rect 8340 16628 8404 16632
rect 9812 16688 9876 16692
rect 9812 16632 9826 16688
rect 9826 16632 9876 16688
rect 9812 16628 9876 16632
rect 9076 16356 9140 16420
rect 11652 16356 11716 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 8892 16220 8956 16284
rect 19748 16084 19812 16148
rect 19380 15812 19444 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 15332 15540 15396 15604
rect 1716 15268 1780 15332
rect 15516 15268 15580 15332
rect 17172 15268 17236 15332
rect 20484 15268 20548 15332
rect 21220 15268 21284 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 7604 15192 7668 15196
rect 7604 15136 7618 15192
rect 7618 15136 7668 15192
rect 7604 15132 7668 15136
rect 24716 15192 24780 15196
rect 24716 15136 24730 15192
rect 24730 15136 24780 15192
rect 24716 15132 24780 15136
rect 12756 14996 12820 15060
rect 1164 14860 1228 14924
rect 17540 14724 17604 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 12756 14588 12820 14652
rect 22140 14588 22204 14652
rect 5580 14180 5644 14244
rect 13860 14180 13924 14244
rect 16436 14240 16500 14244
rect 16436 14184 16450 14240
rect 16450 14184 16500 14240
rect 16436 14180 16500 14184
rect 16620 14180 16684 14244
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 12572 14044 12636 14108
rect 13676 13908 13740 13972
rect 2452 13772 2516 13836
rect 20668 13772 20732 13836
rect 3372 13696 3436 13700
rect 3372 13640 3422 13696
rect 3422 13640 3436 13696
rect 3372 13636 3436 13640
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 5764 13500 5828 13564
rect 17724 13696 17788 13700
rect 17724 13640 17774 13696
rect 17774 13640 17788 13696
rect 17724 13636 17788 13640
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 12388 13500 12452 13564
rect 19380 13560 19444 13564
rect 19380 13504 19394 13560
rect 19394 13504 19444 13560
rect 19380 13500 19444 13504
rect 12204 13228 12268 13292
rect 12388 13228 12452 13292
rect 24532 13288 24596 13292
rect 24532 13232 24582 13288
rect 24582 13232 24596 13288
rect 24532 13228 24596 13232
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 19196 13092 19260 13156
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 22140 13016 22204 13020
rect 22140 12960 22154 13016
rect 22154 12960 22204 13016
rect 22140 12956 22204 12960
rect 4476 12684 4540 12748
rect 3924 12548 3988 12612
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 2084 12336 2148 12340
rect 2084 12280 2134 12336
rect 2134 12280 2148 12336
rect 2084 12276 2148 12280
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 21220 12548 21284 12612
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 12756 11868 12820 11932
rect 15700 11868 15764 11932
rect 20668 11732 20732 11796
rect 8340 11460 8404 11524
rect 15332 11460 15396 11524
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 12756 11324 12820 11388
rect 19748 11324 19812 11388
rect 19012 11052 19076 11116
rect 21036 11052 21100 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 13492 10780 13556 10844
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 14228 10372 14292 10436
rect 19196 10372 19260 10436
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7236 10236 7300 10300
rect 11100 10236 11164 10300
rect 12756 10236 12820 10300
rect 3372 9828 3436 9892
rect 7236 9828 7300 9892
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 980 9692 1044 9756
rect 16620 9692 16684 9756
rect 16988 9616 17052 9620
rect 16988 9560 17002 9616
rect 17002 9560 17052 9616
rect 16988 9556 17052 9560
rect 3372 9420 3436 9484
rect 8524 9284 8588 9348
rect 13860 9284 13924 9348
rect 14596 9284 14660 9348
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 5580 9148 5644 9212
rect 5764 9012 5828 9076
rect 4108 8876 4172 8940
rect 5396 8740 5460 8804
rect 14412 8740 14476 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 7236 8604 7300 8668
rect 2084 8468 2148 8532
rect 14044 8604 14108 8668
rect 15148 8604 15212 8668
rect 15700 8604 15764 8668
rect 2636 8392 2700 8396
rect 2636 8336 2686 8392
rect 2686 8336 2700 8392
rect 2636 8332 2700 8336
rect 12756 8468 12820 8532
rect 14780 8468 14844 8532
rect 12020 8196 12084 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 3372 8060 3436 8124
rect 13676 8060 13740 8124
rect 13860 8060 13924 8124
rect 1348 7924 1412 7988
rect 2452 7984 2516 7988
rect 2452 7928 2466 7984
rect 2466 7928 2516 7984
rect 2452 7924 2516 7928
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 8708 7516 8772 7580
rect 14228 7516 14292 7580
rect 15148 7516 15212 7580
rect 4292 7440 4356 7444
rect 4292 7384 4342 7440
rect 4342 7384 4356 7440
rect 4292 7380 4356 7384
rect 5028 7108 5092 7172
rect 7604 7108 7668 7172
rect 13492 7108 13556 7172
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 12572 6896 12636 6900
rect 12572 6840 12622 6896
rect 12622 6840 12636 6896
rect 12572 6836 12636 6840
rect 5396 6700 5460 6764
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 11100 6428 11164 6492
rect 13492 6488 13556 6492
rect 13492 6432 13542 6488
rect 13542 6432 13556 6488
rect 13492 6428 13556 6432
rect 15516 6488 15580 6492
rect 15516 6432 15530 6488
rect 15530 6432 15580 6488
rect 15516 6428 15580 6432
rect 14964 6020 15028 6084
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 11836 5884 11900 5948
rect 14780 5748 14844 5812
rect 15148 5748 15212 5812
rect 4108 5672 4172 5676
rect 4108 5616 4158 5672
rect 4158 5616 4172 5672
rect 4108 5612 4172 5616
rect 9076 5612 9140 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 12020 5204 12084 5268
rect 3924 4932 3988 4996
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 9812 4796 9876 4860
rect 21220 4856 21284 4860
rect 21220 4800 21234 4856
rect 21234 4800 21284 4856
rect 21220 4796 21284 4800
rect 11836 4660 11900 4724
rect 8524 4448 8588 4452
rect 8524 4392 8538 4448
rect 8538 4392 8588 4448
rect 8524 4388 8588 4392
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 13860 4388 13924 4452
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 1716 4040 1780 4044
rect 1716 3984 1730 4040
rect 1730 3984 1780 4040
rect 1716 3980 1780 3984
rect 3556 3980 3620 4044
rect 5580 3980 5644 4044
rect 17172 4116 17236 4180
rect 19012 3980 19076 4044
rect 20484 3980 20548 4044
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 15332 3708 15396 3772
rect 24532 3708 24596 3772
rect 7788 3572 7852 3636
rect 22324 3572 22388 3636
rect 14964 3436 15028 3500
rect 10916 3300 10980 3364
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 14596 3164 14660 3228
rect 14412 3028 14476 3092
rect 6500 2892 6564 2956
rect 9260 2756 9324 2820
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7236 2620 7300 2684
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 4660 1804 4724 1868
rect 8892 1804 8956 1868
rect 20852 1668 20916 1732
rect 4476 1532 4540 1596
rect 15148 1532 15212 1596
rect 7604 1260 7668 1324
rect 19012 1260 19076 1324
rect 5028 1124 5092 1188
rect 17540 1124 17604 1188
rect 7788 988 7852 1052
rect 16988 988 17052 1052
rect 2636 852 2700 916
rect 1348 716 1412 780
rect 1164 580 1228 644
rect 980 444 1044 508
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 16251 47564 16317 47565
rect 16251 47500 16252 47564
rect 16316 47500 16317 47564
rect 16251 47499 16317 47500
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 15331 42668 15397 42669
rect 15331 42604 15332 42668
rect 15396 42604 15397 42668
rect 15331 42603 15397 42604
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12203 41580 12269 41581
rect 12203 41516 12204 41580
rect 12268 41516 12269 41580
rect 12203 41515 12269 41516
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 11651 25804 11717 25805
rect 11651 25740 11652 25804
rect 11716 25740 11717 25804
rect 11651 25739 11717 25740
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 10915 22540 10981 22541
rect 10915 22476 10916 22540
rect 10980 22476 10981 22540
rect 10915 22475 10981 22476
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 4659 21588 4725 21589
rect 4659 21524 4660 21588
rect 4724 21524 4725 21588
rect 4659 21523 4725 21524
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 3555 18324 3621 18325
rect 3555 18260 3556 18324
rect 3620 18260 3621 18324
rect 3555 18259 3621 18260
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 1715 15332 1781 15333
rect 1715 15268 1716 15332
rect 1780 15268 1781 15332
rect 1715 15267 1781 15268
rect 1163 14924 1229 14925
rect 1163 14860 1164 14924
rect 1228 14860 1229 14924
rect 1163 14859 1229 14860
rect 979 9756 1045 9757
rect 979 9692 980 9756
rect 1044 9692 1045 9756
rect 979 9691 1045 9692
rect 982 509 1042 9691
rect 1166 645 1226 14859
rect 1347 7988 1413 7989
rect 1347 7924 1348 7988
rect 1412 7924 1413 7988
rect 1347 7923 1413 7924
rect 1350 781 1410 7923
rect 1718 4045 1778 15267
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2451 13836 2517 13837
rect 2451 13772 2452 13836
rect 2516 13772 2517 13836
rect 2451 13771 2517 13772
rect 2083 12340 2149 12341
rect 2083 12276 2084 12340
rect 2148 12276 2149 12340
rect 2083 12275 2149 12276
rect 2086 8533 2146 12275
rect 2083 8532 2149 8533
rect 2083 8468 2084 8532
rect 2148 8468 2149 8532
rect 2083 8467 2149 8468
rect 2454 7989 2514 13771
rect 2944 13632 3264 14656
rect 3371 13700 3437 13701
rect 3371 13636 3372 13700
rect 3436 13636 3437 13700
rect 3371 13635 3437 13636
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 3374 9893 3434 13635
rect 3371 9892 3437 9893
rect 3371 9828 3372 9892
rect 3436 9828 3437 9892
rect 3371 9827 3437 9828
rect 3371 9484 3437 9485
rect 3371 9420 3372 9484
rect 3436 9420 3437 9484
rect 3371 9419 3437 9420
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2635 8396 2701 8397
rect 2635 8332 2636 8396
rect 2700 8332 2701 8396
rect 2635 8331 2701 8332
rect 2451 7988 2517 7989
rect 2451 7924 2452 7988
rect 2516 7924 2517 7988
rect 2451 7923 2517 7924
rect 1715 4044 1781 4045
rect 1715 3980 1716 4044
rect 1780 3980 1781 4044
rect 1715 3979 1781 3980
rect 2638 917 2698 8331
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 3374 8125 3434 9419
rect 3371 8124 3437 8125
rect 3371 8060 3372 8124
rect 3436 8060 3437 8124
rect 3371 8059 3437 8060
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 3558 4045 3618 18259
rect 4291 16964 4357 16965
rect 4291 16900 4292 16964
rect 4356 16900 4357 16964
rect 4291 16899 4357 16900
rect 3923 12612 3989 12613
rect 3923 12548 3924 12612
rect 3988 12548 3989 12612
rect 3923 12547 3989 12548
rect 3926 4997 3986 12547
rect 4107 8940 4173 8941
rect 4107 8876 4108 8940
rect 4172 8876 4173 8940
rect 4107 8875 4173 8876
rect 4110 5677 4170 8875
rect 4294 7445 4354 16899
rect 4475 12748 4541 12749
rect 4475 12684 4476 12748
rect 4540 12684 4541 12748
rect 4475 12683 4541 12684
rect 4291 7444 4357 7445
rect 4291 7380 4292 7444
rect 4356 7380 4357 7444
rect 4291 7379 4357 7380
rect 4107 5676 4173 5677
rect 4107 5612 4108 5676
rect 4172 5612 4173 5676
rect 4107 5611 4173 5612
rect 3923 4996 3989 4997
rect 3923 4932 3924 4996
rect 3988 4932 3989 4996
rect 3923 4931 3989 4932
rect 3555 4044 3621 4045
rect 3555 3980 3556 4044
rect 3620 3980 3621 4044
rect 3555 3979 3621 3980
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 4478 1597 4538 12683
rect 4662 1869 4722 21523
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 9259 18052 9325 18053
rect 9259 17988 9260 18052
rect 9324 17988 9325 18052
rect 9259 17987 9325 17988
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 6499 16692 6565 16693
rect 6499 16628 6500 16692
rect 6564 16628 6565 16692
rect 6499 16627 6565 16628
rect 5579 14244 5645 14245
rect 5579 14180 5580 14244
rect 5644 14180 5645 14244
rect 5579 14179 5645 14180
rect 5582 9213 5642 14179
rect 5763 13564 5829 13565
rect 5763 13500 5764 13564
rect 5828 13500 5829 13564
rect 5763 13499 5829 13500
rect 5579 9212 5645 9213
rect 5579 9148 5580 9212
rect 5644 9148 5645 9212
rect 5579 9147 5645 9148
rect 5766 9077 5826 13499
rect 5763 9076 5829 9077
rect 5763 9012 5764 9076
rect 5828 9012 5829 9076
rect 5763 9011 5829 9012
rect 5395 8804 5461 8805
rect 5395 8740 5396 8804
rect 5460 8740 5461 8804
rect 5395 8739 5461 8740
rect 5027 7172 5093 7173
rect 5027 7108 5028 7172
rect 5092 7108 5093 7172
rect 5027 7107 5093 7108
rect 4659 1868 4725 1869
rect 4659 1804 4660 1868
rect 4724 1804 4725 1868
rect 4659 1803 4725 1804
rect 4475 1596 4541 1597
rect 4475 1532 4476 1596
rect 4540 1532 4541 1596
rect 4475 1531 4541 1532
rect 5030 1189 5090 7107
rect 5398 6765 5458 8739
rect 5395 6764 5461 6765
rect 5395 6700 5396 6764
rect 5460 6700 5461 6764
rect 5395 6699 5461 6700
rect 5398 5810 5458 6699
rect 5398 5750 5642 5810
rect 5582 4045 5642 5750
rect 5579 4044 5645 4045
rect 5579 3980 5580 4044
rect 5644 3980 5645 4044
rect 5579 3979 5645 3980
rect 6502 2957 6562 16627
rect 7944 16352 8264 17376
rect 8339 16692 8405 16693
rect 8339 16628 8340 16692
rect 8404 16628 8405 16692
rect 8339 16627 8405 16628
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7603 15196 7669 15197
rect 7603 15132 7604 15196
rect 7668 15132 7669 15196
rect 7603 15131 7669 15132
rect 7235 10300 7301 10301
rect 7235 10236 7236 10300
rect 7300 10236 7301 10300
rect 7235 10235 7301 10236
rect 7238 9893 7298 10235
rect 7235 9892 7301 9893
rect 7235 9828 7236 9892
rect 7300 9828 7301 9892
rect 7235 9827 7301 9828
rect 7235 8668 7301 8669
rect 7235 8604 7236 8668
rect 7300 8604 7301 8668
rect 7235 8603 7301 8604
rect 6499 2956 6565 2957
rect 6499 2892 6500 2956
rect 6564 2892 6565 2956
rect 6499 2891 6565 2892
rect 7238 2685 7298 8603
rect 7606 7173 7666 15131
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 8342 11525 8402 16627
rect 9075 16420 9141 16421
rect 9075 16356 9076 16420
rect 9140 16356 9141 16420
rect 9075 16355 9141 16356
rect 8891 16284 8957 16285
rect 8891 16220 8892 16284
rect 8956 16220 8957 16284
rect 8891 16219 8957 16220
rect 8339 11524 8405 11525
rect 8339 11460 8340 11524
rect 8404 11460 8405 11524
rect 8339 11459 8405 11460
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7603 7172 7669 7173
rect 7603 7108 7604 7172
rect 7668 7108 7669 7172
rect 7603 7107 7669 7108
rect 7235 2684 7301 2685
rect 7235 2620 7236 2684
rect 7300 2620 7301 2684
rect 7235 2619 7301 2620
rect 7606 1325 7666 7107
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7787 3636 7853 3637
rect 7787 3572 7788 3636
rect 7852 3572 7853 3636
rect 7787 3571 7853 3572
rect 7603 1324 7669 1325
rect 7603 1260 7604 1324
rect 7668 1260 7669 1324
rect 7603 1259 7669 1260
rect 5027 1188 5093 1189
rect 5027 1124 5028 1188
rect 5092 1124 5093 1188
rect 5027 1123 5093 1124
rect 7790 1053 7850 3571
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 8342 2790 8402 11459
rect 8894 9690 8954 16219
rect 8710 9630 8954 9690
rect 8523 9348 8589 9349
rect 8523 9284 8524 9348
rect 8588 9284 8589 9348
rect 8523 9283 8589 9284
rect 8526 4453 8586 9283
rect 8710 7581 8770 9630
rect 8707 7580 8773 7581
rect 8707 7516 8708 7580
rect 8772 7516 8773 7580
rect 8707 7515 8773 7516
rect 9078 5677 9138 16355
rect 9075 5676 9141 5677
rect 9075 5612 9076 5676
rect 9140 5612 9141 5676
rect 9075 5611 9141 5612
rect 8523 4452 8589 4453
rect 8523 4388 8524 4452
rect 8588 4388 8589 4452
rect 8523 4387 8589 4388
rect 9262 2821 9322 17987
rect 9811 16692 9877 16693
rect 9811 16628 9812 16692
rect 9876 16628 9877 16692
rect 9811 16627 9877 16628
rect 9814 4861 9874 16627
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 10918 3365 10978 22475
rect 11654 16421 11714 25739
rect 11835 18052 11901 18053
rect 11835 17988 11836 18052
rect 11900 17988 11901 18052
rect 11835 17987 11901 17988
rect 12019 18052 12085 18053
rect 12019 17988 12020 18052
rect 12084 17988 12085 18052
rect 12019 17987 12085 17988
rect 11651 16420 11717 16421
rect 11651 16356 11652 16420
rect 11716 16356 11717 16420
rect 11651 16355 11717 16356
rect 11099 10300 11165 10301
rect 11099 10236 11100 10300
rect 11164 10236 11165 10300
rect 11099 10235 11165 10236
rect 11102 6493 11162 10235
rect 11099 6492 11165 6493
rect 11099 6428 11100 6492
rect 11164 6428 11165 6492
rect 11099 6427 11165 6428
rect 11838 5949 11898 17987
rect 12022 8261 12082 17987
rect 12206 13293 12266 41515
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12571 20908 12637 20909
rect 12571 20844 12572 20908
rect 12636 20844 12637 20908
rect 12571 20843 12637 20844
rect 12574 14109 12634 20843
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12755 15060 12821 15061
rect 12755 14996 12756 15060
rect 12820 14996 12821 15060
rect 12755 14995 12821 14996
rect 12758 14653 12818 14995
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12755 14652 12821 14653
rect 12755 14588 12756 14652
rect 12820 14588 12821 14652
rect 12755 14587 12821 14588
rect 12571 14108 12637 14109
rect 12571 14044 12572 14108
rect 12636 14044 12637 14108
rect 12571 14043 12637 14044
rect 12387 13564 12453 13565
rect 12387 13500 12388 13564
rect 12452 13500 12453 13564
rect 12387 13499 12453 13500
rect 12390 13293 12450 13499
rect 12203 13292 12269 13293
rect 12203 13228 12204 13292
rect 12268 13228 12269 13292
rect 12203 13227 12269 13228
rect 12387 13292 12453 13293
rect 12387 13228 12388 13292
rect 12452 13228 12453 13292
rect 12387 13227 12453 13228
rect 12019 8260 12085 8261
rect 12019 8196 12020 8260
rect 12084 8196 12085 8260
rect 12019 8195 12085 8196
rect 11835 5948 11901 5949
rect 11835 5884 11836 5948
rect 11900 5884 11901 5948
rect 11835 5883 11901 5884
rect 11838 4725 11898 5883
rect 12022 5269 12082 8195
rect 12574 6901 12634 14043
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12755 11932 12821 11933
rect 12755 11868 12756 11932
rect 12820 11868 12821 11932
rect 12755 11867 12821 11868
rect 12758 11389 12818 11867
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12755 11388 12821 11389
rect 12755 11324 12756 11388
rect 12820 11324 12821 11388
rect 12755 11323 12821 11324
rect 12944 10368 13264 11392
rect 13494 10845 13554 23427
rect 14227 20772 14293 20773
rect 14227 20708 14228 20772
rect 14292 20708 14293 20772
rect 14227 20707 14293 20708
rect 14043 18052 14109 18053
rect 14043 17988 14044 18052
rect 14108 17988 14109 18052
rect 14043 17987 14109 17988
rect 13859 14244 13925 14245
rect 13859 14180 13860 14244
rect 13924 14180 13925 14244
rect 13859 14179 13925 14180
rect 13675 13972 13741 13973
rect 13675 13908 13676 13972
rect 13740 13908 13741 13972
rect 13675 13907 13741 13908
rect 13491 10844 13557 10845
rect 13491 10780 13492 10844
rect 13556 10780 13557 10844
rect 13491 10779 13557 10780
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12755 10300 12821 10301
rect 12755 10236 12756 10300
rect 12820 10236 12821 10300
rect 12755 10235 12821 10236
rect 12758 8533 12818 10235
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12755 8532 12821 8533
rect 12755 8468 12756 8532
rect 12820 8468 12821 8532
rect 12755 8467 12821 8468
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 13494 7173 13554 10779
rect 13678 8125 13738 13907
rect 13862 9349 13922 14179
rect 13859 9348 13925 9349
rect 13859 9284 13860 9348
rect 13924 9284 13925 9348
rect 13859 9283 13925 9284
rect 14046 8669 14106 17987
rect 14230 12450 14290 20707
rect 14963 19684 15029 19685
rect 14963 19620 14964 19684
rect 15028 19620 15029 19684
rect 14963 19619 15029 19620
rect 14966 19005 15026 19619
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 14963 19004 15029 19005
rect 14963 18940 14964 19004
rect 15028 18940 15029 19004
rect 14963 18939 15029 18940
rect 15150 18869 15210 19347
rect 15147 18868 15213 18869
rect 15147 18804 15148 18868
rect 15212 18804 15213 18868
rect 15147 18803 15213 18804
rect 15334 15605 15394 42603
rect 15699 34508 15765 34509
rect 15699 34444 15700 34508
rect 15764 34444 15765 34508
rect 15699 34443 15765 34444
rect 15702 17917 15762 34443
rect 16254 25397 16314 47499
rect 17944 46816 18264 47840
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 21035 47700 21101 47701
rect 21035 47636 21036 47700
rect 21100 47636 21101 47700
rect 21035 47635 21101 47636
rect 20483 47020 20549 47021
rect 20483 46956 20484 47020
rect 20548 46956 20549 47020
rect 20483 46955 20549 46956
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 19747 40084 19813 40085
rect 19747 40020 19748 40084
rect 19812 40020 19813 40084
rect 19747 40019 19813 40020
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 16435 35868 16501 35869
rect 16435 35804 16436 35868
rect 16500 35804 16501 35868
rect 16435 35803 16501 35804
rect 16251 25396 16317 25397
rect 16251 25332 16252 25396
rect 16316 25332 16317 25396
rect 16251 25331 16317 25332
rect 15883 18052 15949 18053
rect 15883 17988 15884 18052
rect 15948 17988 15949 18052
rect 15883 17987 15949 17988
rect 15699 17916 15765 17917
rect 15699 17852 15700 17916
rect 15764 17852 15765 17916
rect 15699 17851 15765 17852
rect 15886 16010 15946 17987
rect 15702 15950 15946 16010
rect 15331 15604 15397 15605
rect 15331 15540 15332 15604
rect 15396 15540 15397 15604
rect 15331 15539 15397 15540
rect 15515 15332 15581 15333
rect 15515 15268 15516 15332
rect 15580 15268 15581 15332
rect 15515 15267 15581 15268
rect 14230 12390 14474 12450
rect 14227 10436 14293 10437
rect 14227 10372 14228 10436
rect 14292 10372 14293 10436
rect 14227 10371 14293 10372
rect 14043 8668 14109 8669
rect 14043 8604 14044 8668
rect 14108 8604 14109 8668
rect 14043 8603 14109 8604
rect 13675 8124 13741 8125
rect 13675 8060 13676 8124
rect 13740 8060 13741 8124
rect 13675 8059 13741 8060
rect 13859 8124 13925 8125
rect 13859 8060 13860 8124
rect 13924 8060 13925 8124
rect 13859 8059 13925 8060
rect 13491 7172 13557 7173
rect 13491 7108 13492 7172
rect 13556 7108 13557 7172
rect 13491 7107 13557 7108
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12571 6900 12637 6901
rect 12571 6836 12572 6900
rect 12636 6836 12637 6900
rect 12571 6835 12637 6836
rect 12944 6016 13264 7040
rect 13494 6493 13554 7107
rect 13491 6492 13557 6493
rect 13491 6428 13492 6492
rect 13556 6428 13557 6492
rect 13491 6427 13557 6428
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12019 5268 12085 5269
rect 12019 5204 12020 5268
rect 12084 5204 12085 5268
rect 12019 5203 12085 5204
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 11835 4724 11901 4725
rect 11835 4660 11836 4724
rect 11900 4660 11901 4724
rect 11835 4659 11901 4660
rect 12944 3840 13264 4864
rect 13862 4453 13922 8059
rect 14230 7581 14290 10371
rect 14414 8805 14474 12390
rect 15331 11524 15397 11525
rect 15331 11460 15332 11524
rect 15396 11460 15397 11524
rect 15331 11459 15397 11460
rect 14595 9348 14661 9349
rect 14595 9284 14596 9348
rect 14660 9284 14661 9348
rect 14595 9283 14661 9284
rect 14411 8804 14477 8805
rect 14411 8740 14412 8804
rect 14476 8740 14477 8804
rect 14411 8739 14477 8740
rect 14227 7580 14293 7581
rect 14227 7516 14228 7580
rect 14292 7516 14293 7580
rect 14227 7515 14293 7516
rect 13859 4452 13925 4453
rect 13859 4388 13860 4452
rect 13924 4388 13925 4452
rect 13859 4387 13925 4388
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 10915 3364 10981 3365
rect 10915 3300 10916 3364
rect 10980 3300 10981 3364
rect 10915 3299 10981 3300
rect 9259 2820 9325 2821
rect 8342 2730 8954 2790
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 8894 1869 8954 2730
rect 12944 2752 13264 3776
rect 14414 3093 14474 8739
rect 14598 3229 14658 9283
rect 15147 8668 15213 8669
rect 15147 8604 15148 8668
rect 15212 8604 15213 8668
rect 15147 8603 15213 8604
rect 14779 8532 14845 8533
rect 14779 8468 14780 8532
rect 14844 8468 14845 8532
rect 14779 8467 14845 8468
rect 14782 5813 14842 8467
rect 15150 7581 15210 8603
rect 15147 7580 15213 7581
rect 15147 7516 15148 7580
rect 15212 7516 15213 7580
rect 15147 7515 15213 7516
rect 14963 6084 15029 6085
rect 14963 6020 14964 6084
rect 15028 6020 15029 6084
rect 14963 6019 15029 6020
rect 14779 5812 14845 5813
rect 14779 5748 14780 5812
rect 14844 5748 14845 5812
rect 14779 5747 14845 5748
rect 14966 3501 15026 6019
rect 15147 5812 15213 5813
rect 15147 5748 15148 5812
rect 15212 5748 15213 5812
rect 15147 5747 15213 5748
rect 14963 3500 15029 3501
rect 14963 3436 14964 3500
rect 15028 3436 15029 3500
rect 14963 3435 15029 3436
rect 14595 3228 14661 3229
rect 14595 3164 14596 3228
rect 14660 3164 14661 3228
rect 14595 3163 14661 3164
rect 14411 3092 14477 3093
rect 14411 3028 14412 3092
rect 14476 3028 14477 3092
rect 14411 3027 14477 3028
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 8891 1868 8957 1869
rect 8891 1804 8892 1868
rect 8956 1804 8957 1868
rect 8891 1803 8957 1804
rect 15150 1597 15210 5747
rect 15334 3773 15394 11459
rect 15518 6493 15578 15267
rect 15702 11933 15762 15950
rect 16438 14245 16498 35803
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 18643 30836 18709 30837
rect 18643 30772 18644 30836
rect 18708 30772 18709 30836
rect 18643 30771 18709 30772
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 18646 27573 18706 30771
rect 18643 27572 18709 27573
rect 18643 27508 18644 27572
rect 18708 27508 18709 27572
rect 18643 27507 18709 27508
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17723 26484 17789 26485
rect 17723 26420 17724 26484
rect 17788 26420 17789 26484
rect 17723 26419 17789 26420
rect 17539 21180 17605 21181
rect 17539 21116 17540 21180
rect 17604 21116 17605 21180
rect 17539 21115 17605 21116
rect 16987 19140 17053 19141
rect 16987 19076 16988 19140
rect 17052 19076 17053 19140
rect 16987 19075 17053 19076
rect 16435 14244 16501 14245
rect 16435 14180 16436 14244
rect 16500 14180 16501 14244
rect 16435 14179 16501 14180
rect 16619 14244 16685 14245
rect 16619 14180 16620 14244
rect 16684 14180 16685 14244
rect 16619 14179 16685 14180
rect 15699 11932 15765 11933
rect 15699 11868 15700 11932
rect 15764 11868 15765 11932
rect 15699 11867 15765 11868
rect 15702 8669 15762 11867
rect 16622 9757 16682 14179
rect 16619 9756 16685 9757
rect 16619 9692 16620 9756
rect 16684 9692 16685 9756
rect 16619 9691 16685 9692
rect 16990 9621 17050 19075
rect 17171 15332 17237 15333
rect 17171 15268 17172 15332
rect 17236 15268 17237 15332
rect 17171 15267 17237 15268
rect 16987 9620 17053 9621
rect 16987 9556 16988 9620
rect 17052 9556 17053 9620
rect 16987 9555 17053 9556
rect 15699 8668 15765 8669
rect 15699 8604 15700 8668
rect 15764 8604 15765 8668
rect 15699 8603 15765 8604
rect 15515 6492 15581 6493
rect 15515 6428 15516 6492
rect 15580 6428 15581 6492
rect 15515 6427 15581 6428
rect 17174 4181 17234 15267
rect 17542 14789 17602 21115
rect 17539 14788 17605 14789
rect 17539 14724 17540 14788
rect 17604 14724 17605 14788
rect 17539 14723 17605 14724
rect 17726 13701 17786 26419
rect 17944 26144 18264 27168
rect 19011 26348 19077 26349
rect 19011 26284 19012 26348
rect 19076 26284 19077 26348
rect 19011 26283 19077 26284
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17723 13700 17789 13701
rect 17723 13636 17724 13700
rect 17788 13636 17789 13700
rect 17723 13635 17789 13636
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 19014 11117 19074 26283
rect 19750 16149 19810 40019
rect 20486 21453 20546 46955
rect 21038 25397 21098 47635
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22691 29068 22757 29069
rect 22691 29004 22692 29068
rect 22756 29004 22757 29068
rect 22691 29003 22757 29004
rect 21035 25396 21101 25397
rect 21035 25332 21036 25396
rect 21100 25332 21101 25396
rect 21035 25331 21101 25332
rect 20851 24988 20917 24989
rect 20851 24924 20852 24988
rect 20916 24924 20917 24988
rect 20851 24923 20917 24924
rect 22139 24988 22205 24989
rect 22139 24924 22140 24988
rect 22204 24924 22205 24988
rect 22139 24923 22205 24924
rect 20483 21452 20549 21453
rect 20483 21388 20484 21452
rect 20548 21388 20549 21452
rect 20483 21387 20549 21388
rect 19747 16148 19813 16149
rect 19747 16084 19748 16148
rect 19812 16084 19813 16148
rect 19747 16083 19813 16084
rect 19379 15876 19445 15877
rect 19379 15812 19380 15876
rect 19444 15812 19445 15876
rect 19379 15811 19445 15812
rect 19382 13565 19442 15811
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19195 13156 19261 13157
rect 19195 13092 19196 13156
rect 19260 13092 19261 13156
rect 19195 13091 19261 13092
rect 19011 11116 19077 11117
rect 19011 11052 19012 11116
rect 19076 11052 19077 11116
rect 19011 11051 19077 11052
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 19198 10437 19258 13091
rect 19750 11389 19810 16083
rect 20486 15333 20546 21387
rect 20667 19684 20733 19685
rect 20667 19620 20668 19684
rect 20732 19620 20733 19684
rect 20667 19619 20733 19620
rect 20483 15332 20549 15333
rect 20483 15268 20484 15332
rect 20548 15268 20549 15332
rect 20483 15267 20549 15268
rect 20670 14650 20730 19619
rect 20486 14590 20730 14650
rect 19747 11388 19813 11389
rect 19747 11324 19748 11388
rect 19812 11324 19813 11388
rect 19747 11323 19813 11324
rect 19195 10436 19261 10437
rect 19195 10372 19196 10436
rect 19260 10372 19261 10436
rect 19195 10371 19261 10372
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17171 4180 17237 4181
rect 17171 4116 17172 4180
rect 17236 4116 17237 4180
rect 17171 4115 17237 4116
rect 15331 3772 15397 3773
rect 15331 3708 15332 3772
rect 15396 3708 15397 3772
rect 15331 3707 15397 3708
rect 17944 3296 18264 4320
rect 20486 4045 20546 14590
rect 20667 13836 20733 13837
rect 20667 13772 20668 13836
rect 20732 13772 20733 13836
rect 20667 13771 20733 13772
rect 20670 11797 20730 13771
rect 20667 11796 20733 11797
rect 20667 11732 20668 11796
rect 20732 11732 20733 11796
rect 20667 11731 20733 11732
rect 19011 4044 19077 4045
rect 19011 3980 19012 4044
rect 19076 3980 19077 4044
rect 19011 3979 19077 3980
rect 20483 4044 20549 4045
rect 20483 3980 20484 4044
rect 20548 3980 20549 4044
rect 20483 3979 20549 3980
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 15147 1596 15213 1597
rect 15147 1532 15148 1596
rect 15212 1532 15213 1596
rect 15147 1531 15213 1532
rect 19014 1325 19074 3979
rect 20854 1733 20914 24923
rect 21035 19004 21101 19005
rect 21035 18940 21036 19004
rect 21100 18940 21101 19004
rect 21035 18939 21101 18940
rect 21038 11117 21098 18939
rect 21219 15332 21285 15333
rect 21219 15268 21220 15332
rect 21284 15268 21285 15332
rect 21219 15267 21285 15268
rect 21222 12613 21282 15267
rect 22142 14653 22202 24923
rect 22323 17916 22389 17917
rect 22323 17852 22324 17916
rect 22388 17852 22389 17916
rect 22323 17851 22389 17852
rect 22139 14652 22205 14653
rect 22139 14588 22140 14652
rect 22204 14588 22205 14652
rect 22139 14587 22205 14588
rect 22142 13021 22202 14587
rect 22139 13020 22205 13021
rect 22139 12956 22140 13020
rect 22204 12956 22205 13020
rect 22139 12955 22205 12956
rect 21219 12612 21285 12613
rect 21219 12548 21220 12612
rect 21284 12548 21285 12612
rect 21219 12547 21285 12548
rect 21035 11116 21101 11117
rect 21035 11052 21036 11116
rect 21100 11052 21101 11116
rect 21035 11051 21101 11052
rect 21222 4861 21282 12547
rect 21219 4860 21285 4861
rect 21219 4796 21220 4860
rect 21284 4796 21285 4860
rect 21219 4795 21285 4796
rect 22326 3637 22386 17851
rect 22694 17373 22754 29003
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 24715 25396 24781 25397
rect 24715 25332 24716 25396
rect 24780 25332 24781 25396
rect 24715 25331 24781 25332
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 24531 22676 24597 22677
rect 24531 22612 24532 22676
rect 24596 22612 24597 22676
rect 24531 22611 24597 22612
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22691 17372 22757 17373
rect 22691 17308 22692 17372
rect 22756 17308 22757 17372
rect 22691 17307 22757 17308
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 24534 13293 24594 22611
rect 24718 15197 24778 25331
rect 24715 15196 24781 15197
rect 24715 15132 24716 15196
rect 24780 15132 24781 15196
rect 24715 15131 24781 15132
rect 24531 13292 24597 13293
rect 24531 13228 24532 13292
rect 24596 13228 24597 13292
rect 24531 13227 24597 13228
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22323 3636 22389 3637
rect 22323 3572 22324 3636
rect 22388 3572 22389 3636
rect 22323 3571 22389 3572
rect 22944 2752 23264 3776
rect 24534 3773 24594 13227
rect 24531 3772 24597 3773
rect 24531 3708 24532 3772
rect 24596 3708 24597 3772
rect 24531 3707 24597 3708
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 20851 1732 20917 1733
rect 20851 1668 20852 1732
rect 20916 1668 20917 1732
rect 20851 1667 20917 1668
rect 19011 1324 19077 1325
rect 19011 1260 19012 1324
rect 19076 1260 19077 1324
rect 19011 1259 19077 1260
rect 17539 1188 17605 1189
rect 17539 1124 17540 1188
rect 17604 1124 17605 1188
rect 17539 1123 17605 1124
rect 7787 1052 7853 1053
rect 7787 988 7788 1052
rect 7852 988 7853 1052
rect 7787 987 7853 988
rect 16987 1052 17053 1053
rect 16987 988 16988 1052
rect 17052 1050 17053 1052
rect 17542 1050 17602 1123
rect 17052 990 17602 1050
rect 17052 988 17053 990
rect 16987 987 17053 988
rect 2635 916 2701 917
rect 2635 852 2636 916
rect 2700 852 2701 916
rect 2635 851 2701 852
rect 1347 780 1413 781
rect 1347 716 1348 780
rect 1412 716 1413 780
rect 1347 715 1413 716
rect 1163 644 1229 645
rect 1163 580 1164 644
rect 1228 580 1229 644
rect 1163 579 1229 580
rect 979 508 1045 509
rect 979 444 980 508
rect 1044 444 1045 508
rect 979 443 1045 444
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3496 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1679235063
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1679235063
transform 1 0 3864 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1679235063
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform 1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1679235063
transform 1 0 14720 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1679235063
transform 1 0 3128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 3128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform 1 0 2944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 3956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _123_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1679235063
transform 1 0 3680 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1679235063
transform 1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1679235063
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1679235063
transform 1 0 5980 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1679235063
transform 1 0 21804 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform 1 0 21068 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 21988 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 20976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 20608 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 18492 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 16008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 6624 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1679235063
transform 1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1679235063
transform 1 0 3128 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1679235063
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1679235063
transform 1 0 14260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1679235063
transform 1 0 4968 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 6532 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1679235063
transform 1 0 7636 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1679235063
transform 1 0 8648 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 7084 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 9016 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1679235063
transform 1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1679235063
transform 1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1679235063
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1679235063
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1679235063
transform 1 0 13064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1679235063
transform 1 0 7084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1679235063
transform 1 0 22080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1679235063
transform 1 0 20240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1679235063
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1679235063
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1679235063
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1679235063
transform 1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform 1 0 25208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1679235063
transform 1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1679235063
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1679235063
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform 1 0 23276 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 14168 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1679235063
transform 1 0 11592 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1679235063
transform 1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 15640 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 2392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1679235063
transform 1 0 2024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1679235063
transform 1 0 1932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1679235063
transform 1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1679235063
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1679235063
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 10672 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 18860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 17296 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 15364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 9384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16008 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 12512 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 11040 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11868 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 10856 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 11132 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 8280 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 8556 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8280 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 20424 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 16192 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 15548 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 16836 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 23184 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 23368 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 21436 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout143_A
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout144_A
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout145_A
timestamp 1679235063
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout146_A
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout147_A
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout148_A
timestamp 1679235063
transform 1 0 20700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout149_A
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout151_A
timestamp 1679235063
transform 1 0 21160 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout152_A
timestamp 1679235063
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout153_A
timestamp 1679235063
transform 1 0 23460 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold29_A
timestamp 1679235063
transform 1 0 9016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold46_A
timestamp 1679235063
transform 1 0 9016 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold65_A
timestamp 1679235063
transform 1 0 1472 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold104_A
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold170_A
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold243_A
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold244_A
timestamp 1679235063
transform 1 0 4968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold245_A
timestamp 1679235063
transform 1 0 6440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold246_A
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold249_A
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold250_A
timestamp 1679235063
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold253_A
timestamp 1679235063
transform 1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold259_A
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold260_A
timestamp 1679235063
transform 1 0 3864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold265_A
timestamp 1679235063
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold285_A
timestamp 1679235063
transform 1 0 5704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold287_A
timestamp 1679235063
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold304_A
timestamp 1679235063
transform 1 0 16928 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold305_A
timestamp 1679235063
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold314_A
timestamp 1679235063
transform 1 0 16192 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold318_A
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold327_A
timestamp 1679235063
transform 1 0 1472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold338_A
timestamp 1679235063
transform 1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold343_A
timestamp 1679235063
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 23460 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 24932 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 24748 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 24564 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 24656 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 24104 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 24656 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 12052 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 24656 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 24656 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 24748 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 24748 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 24656 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 16008 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 23736 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 18492 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 18124 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 1656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 1472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 2024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 1472 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 3680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 1472 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 2392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 2576 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 6440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 1840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 1472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 2944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 1472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 1472 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 1564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 1472 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 6256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 15364 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 17296 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 18124 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 24472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 23920 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 23736 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 24472 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 22356 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 21988 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 24104 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1679235063
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1679235063
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1679235063
transform 1 0 23644 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1679235063
transform 1 0 17848 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1679235063
transform 1 0 23736 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output85_A
timestamp 1679235063
transform 1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1679235063
transform 1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1679235063
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1679235063
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output104_A
timestamp 1679235063
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output105_A
timestamp 1679235063
transform 1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output106_A
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1679235063
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1679235063
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1679235063
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1679235063
transform 1 0 1472 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1679235063
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1679235063
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1679235063
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1679235063
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 23460 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23000 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22540 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11868 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11592 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13064 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16008 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15088 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15732 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16008 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 24012 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 23828 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 1472 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 20056 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 2208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21988 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24104 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23552 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20516 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20332 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21620 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4784 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23920 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4968 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21712 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 13524 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20516 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23736 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16192 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 18860 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18676 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 18860 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16284 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 10580 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19044 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16652 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16744 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11500 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18860 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 10580 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14352 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 14260 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 10120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16100 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17848 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18032 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17480 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17664 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16284 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17020 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22264 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 21068 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 21160 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23184 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 23000 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 25024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 21620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 17848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9108 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6716 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6348 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7912 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9292 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6624 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8004 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10120 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8004 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8188 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 8648 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13984 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14536 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 11776 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11316 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__197 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9752 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9292 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14720 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15272 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12788 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12696 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9752 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10212 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__198
timestamp 1679235063
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9200 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 8648 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9016 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12052 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__199
timestamp 1679235063
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14720 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10396 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9108 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14444 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 13248 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12696 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11776 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 15640 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__200
timestamp 1679235063
transform 1 0 15824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10028 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9660 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15548 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13248 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11684 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 10580 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 14444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 12420 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 10212 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 9292 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9660 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 14260 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 11408 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 10028 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 8648 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 12144 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 10212 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 7452 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 7728 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15916 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 12512 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 10488 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 12420 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 18032 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 19596 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 17756 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 19688 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 14260 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 14812 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 14352 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 15364 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 20792 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21896 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 19872 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout143 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout144
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout145 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout146
timestamp 1679235063
transform 1 0 12788 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout147
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout148
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout149
timestamp 1679235063
transform 1 0 22080 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout150
timestamp 1679235063
transform 1 0 19412 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout151 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18400 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout152
timestamp 1679235063
transform 1 0 20976 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout153
timestamp 1679235063
transform 1 0 22080 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1679235063
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43
timestamp 1679235063
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1679235063
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1679235063
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1679235063
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_165
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_243
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1679235063
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1679235063
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1679235063
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1679235063
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_51
timestamp 1679235063
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1679235063
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1679235063
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1679235063
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1679235063
transform 1 0 10120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1679235063
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1679235063
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1679235063
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1679235063
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_263
timestamp 1679235063
transform 1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1679235063
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1679235063
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1679235063
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1679235063
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1679235063
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1679235063
transform 1 0 10488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_114
timestamp 1679235063
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_120
timestamp 1679235063
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1679235063
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1679235063
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1679235063
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1679235063
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_239
timestamp 1679235063
transform 1 0 23092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_249
timestamp 1679235063
transform 1 0 24012 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_264
timestamp 1679235063
transform 1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1679235063
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1679235063
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_48
timestamp 1679235063
transform 1 0 5520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1679235063
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1679235063
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1679235063
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1679235063
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1679235063
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_115
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1679235063
transform 1 0 11960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1679235063
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_160
timestamp 1679235063
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_171
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_182
timestamp 1679235063
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_206
timestamp 1679235063
transform 1 0 20056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1679235063
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1679235063
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1679235063
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_20
timestamp 1679235063
transform 1 0 2944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1679235063
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1679235063
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1679235063
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1679235063
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1679235063
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1679235063
transform 1 0 10488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1679235063
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_126
timestamp 1679235063
transform 1 0 12696 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1679235063
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1679235063
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1679235063
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1679235063
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_205
timestamp 1679235063
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1679235063
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_263
timestamp 1679235063
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1679235063
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_25
timestamp 1679235063
transform 1 0 3404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_29
timestamp 1679235063
transform 1 0 3772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1679235063
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1679235063
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1679235063
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1679235063
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1679235063
transform 1 0 7912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1679235063
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1679235063
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1679235063
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_115
timestamp 1679235063
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1679235063
transform 1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_150
timestamp 1679235063
transform 1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1679235063
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1679235063
transform 1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1679235063
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1679235063
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_217
timestamp 1679235063
transform 1 0 21068 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1679235063
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1679235063
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1679235063
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1679235063
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1679235063
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_39
timestamp 1679235063
transform 1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1679235063
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1679235063
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1679235063
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1679235063
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1679235063
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 1679235063
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1679235063
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_123
timestamp 1679235063
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp 1679235063
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1679235063
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1679235063
transform 1 0 14536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1679235063
transform 1 0 15640 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1679235063
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1679235063
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1679235063
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_239
timestamp 1679235063
transform 1 0 23092 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_264
timestamp 1679235063
transform 1 0 25392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1679235063
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1679235063
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_32
timestamp 1679235063
transform 1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1679235063
transform 1 0 4416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1679235063
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1679235063
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1679235063
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1679235063
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1679235063
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1679235063
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1679235063
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1679235063
transform 1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_180
timestamp 1679235063
transform 1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1679235063
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1679235063
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_219
timestamp 1679235063
transform 1 0 21252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1679235063
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1679235063
transform 1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1679235063
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1679235063
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1679235063
transform 1 0 4692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1679235063
transform 1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1679235063
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1679235063
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1679235063
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_89
timestamp 1679235063
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1679235063
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_123
timestamp 1679235063
transform 1 0 12420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1679235063
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1679235063
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1679235063
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1679235063
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_164
timestamp 1679235063
transform 1 0 16192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_174
timestamp 1679235063
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1679235063
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1679235063
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1679235063
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1679235063
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1679235063
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1679235063
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1679235063
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 1679235063
transform 1 0 4968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1679235063
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_61
timestamp 1679235063
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1679235063
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1679235063
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp 1679235063
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_130
timestamp 1679235063
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1679235063
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1679235063
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1679235063
transform 1 0 17112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_180
timestamp 1679235063
transform 1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1679235063
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_247
timestamp 1679235063
transform 1 0 23828 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_263
timestamp 1679235063
transform 1 0 25300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_5
timestamp 1679235063
transform 1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1679235063
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1679235063
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1679235063
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1679235063
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1679235063
transform 1 0 4968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1679235063
transform 1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_58
timestamp 1679235063
transform 1 0 6440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1679235063
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1679235063
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1679235063
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 1679235063
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1679235063
transform 1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_131
timestamp 1679235063
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1679235063
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_156
timestamp 1679235063
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1679235063
transform 1 0 16468 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1679235063
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 1679235063
transform 1 0 20240 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1679235063
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1679235063
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_263
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_5
timestamp 1679235063
transform 1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1679235063
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1679235063
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1679235063
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1679235063
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1679235063
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1679235063
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1679235063
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1679235063
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1679235063
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1679235063
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp 1679235063
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1679235063
transform 1 0 15364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_180
timestamp 1679235063
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1679235063
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1679235063
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1679235063
transform 1 0 1656 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1679235063
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_18
timestamp 1679235063
transform 1 0 2760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1679235063
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1679235063
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1679235063
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1679235063
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1679235063
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1679235063
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1679235063
transform 1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1679235063
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_116
timestamp 1679235063
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1679235063
transform 1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_143
timestamp 1679235063
transform 1 0 14260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_146
timestamp 1679235063
transform 1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1679235063
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1679235063
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_201
timestamp 1679235063
transform 1 0 19596 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1679235063
transform 1 0 21712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1679235063
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_12
timestamp 1679235063
transform 1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1679235063
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_26
timestamp 1679235063
transform 1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1679235063
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1679235063
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1679235063
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_68
timestamp 1679235063
transform 1 0 7360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_80
timestamp 1679235063
transform 1 0 8464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1679235063
transform 1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1679235063
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_142
timestamp 1679235063
transform 1 0 14168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1679235063
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_159
timestamp 1679235063
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1679235063
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1679235063
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1679235063
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_190
timestamp 1679235063
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_202
timestamp 1679235063
transform 1 0 19688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1679235063
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_21
timestamp 1679235063
transform 1 0 3036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1679235063
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1679235063
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1679235063
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1679235063
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1679235063
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1679235063
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_108
timestamp 1679235063
transform 1 0 11040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_114
timestamp 1679235063
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1679235063
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1679235063
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_171
timestamp 1679235063
transform 1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_182
timestamp 1679235063
transform 1 0 17848 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1679235063
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_211
timestamp 1679235063
transform 1 0 20516 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_232
timestamp 1679235063
transform 1 0 22448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_245
timestamp 1679235063
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1679235063
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_263
timestamp 1679235063
transform 1 0 25300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1679235063
transform 1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1679235063
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1679235063
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1679235063
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1679235063
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1679235063
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1679235063
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1679235063
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_70
timestamp 1679235063
transform 1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1679235063
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1679235063
transform 1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1679235063
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1679235063
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1679235063
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_148
timestamp 1679235063
transform 1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1679235063
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_171
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1679235063
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1679235063
transform 1 0 18952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_198
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_234
timestamp 1679235063
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_258
timestamp 1679235063
transform 1 0 24840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_8
timestamp 1679235063
transform 1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_14
timestamp 1679235063
transform 1 0 2392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1679235063
transform 1 0 2852 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1679235063
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1679235063
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_42
timestamp 1679235063
transform 1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1679235063
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1679235063
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1679235063
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_95
timestamp 1679235063
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_108
timestamp 1679235063
transform 1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1679235063
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1679235063
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1679235063
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1679235063
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1679235063
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_175
timestamp 1679235063
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_180
timestamp 1679235063
transform 1 0 17664 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1679235063
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1679235063
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_222
timestamp 1679235063
transform 1 0 21528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1679235063
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_6
timestamp 1679235063
transform 1 0 1656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1679235063
transform 1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_18
timestamp 1679235063
transform 1 0 2760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1679235063
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1679235063
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1679235063
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1679235063
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1679235063
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1679235063
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1679235063
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1679235063
transform 1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1679235063
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1679235063
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_154
timestamp 1679235063
transform 1 0 15272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1679235063
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_195
timestamp 1679235063
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1679235063
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1679235063
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1679235063
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1679235063
transform 1 0 1748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_12
timestamp 1679235063
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_19
timestamp 1679235063
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1679235063
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_34
timestamp 1679235063
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_46
timestamp 1679235063
transform 1 0 5336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1679235063
transform 1 0 6440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1679235063
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1679235063
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1679235063
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1679235063
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1679235063
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_135
timestamp 1679235063
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1679235063
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1679235063
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1679235063
transform 1 0 16744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_182
timestamp 1679235063
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1679235063
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1679235063
transform 1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_231
timestamp 1679235063
transform 1 0 22356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_243
timestamp 1679235063
transform 1 0 23460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_263
timestamp 1679235063
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1679235063
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1679235063
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_19
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1679235063
transform 1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1679235063
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_42
timestamp 1679235063
transform 1 0 4968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1679235063
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_63
timestamp 1679235063
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1679235063
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1679235063
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1679235063
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1679235063
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_143
timestamp 1679235063
transform 1 0 14260 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1679235063
transform 1 0 18676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1679235063
transform 1 0 19412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_212
timestamp 1679235063
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_220
timestamp 1679235063
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1679235063
transform 1 0 22632 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1679235063
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_8
timestamp 1679235063
transform 1 0 1840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1679235063
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_24
timestamp 1679235063
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_35
timestamp 1679235063
transform 1 0 4324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1679235063
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1679235063
transform 1 0 6348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1679235063
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1679235063
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1679235063
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 1679235063
transform 1 0 10304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1679235063
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1679235063
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1679235063
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1679235063
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1679235063
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1679235063
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_182
timestamp 1679235063
transform 1 0 17848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1679235063
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1679235063
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1679235063
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_263
timestamp 1679235063
transform 1 0 25300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1679235063
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1679235063
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1679235063
transform 1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1679235063
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1679235063
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_81
timestamp 1679235063
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1679235063
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1679235063
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1679235063
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1679235063
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1679235063
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_180
timestamp 1679235063
transform 1 0 17664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_186
timestamp 1679235063
transform 1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1679235063
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1679235063
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1679235063
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_231
timestamp 1679235063
transform 1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1679235063
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_263
timestamp 1679235063
transform 1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1679235063
transform 1 0 1656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1679235063
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_19
timestamp 1679235063
transform 1 0 2852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1679235063
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1679235063
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1679235063
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1679235063
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_89
timestamp 1679235063
transform 1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_94
timestamp 1679235063
transform 1 0 9752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_121
timestamp 1679235063
transform 1 0 12236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1679235063
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_153
timestamp 1679235063
transform 1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_159
timestamp 1679235063
transform 1 0 15732 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_169
timestamp 1679235063
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1679235063
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_185
timestamp 1679235063
transform 1 0 18124 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_208
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1679235063
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_227
timestamp 1679235063
transform 1 0 21988 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_263
timestamp 1679235063
transform 1 0 25300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_13
timestamp 1679235063
transform 1 0 2300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_20
timestamp 1679235063
transform 1 0 2944 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1679235063
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1679235063
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_61
timestamp 1679235063
transform 1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1679235063
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1679235063
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1679235063
transform 1 0 12420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1679235063
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_151
timestamp 1679235063
transform 1 0 14996 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1679235063
transform 1 0 15456 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 1679235063
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1679235063
transform 1 0 18032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1679235063
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1679235063
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1679235063
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_251
timestamp 1679235063
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_263
timestamp 1679235063
transform 1 0 25300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_34
timestamp 1679235063
transform 1 0 4232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1679235063
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1679235063
transform 1 0 6256 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_80
timestamp 1679235063
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1679235063
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_103
timestamp 1679235063
transform 1 0 10580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_107
timestamp 1679235063
transform 1 0 10948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1679235063
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1679235063
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1679235063
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_160
timestamp 1679235063
transform 1 0 15824 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_164
timestamp 1679235063
transform 1 0 16192 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1679235063
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1679235063
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1679235063
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 1679235063
transform 1 0 20148 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_264
timestamp 1679235063
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1656 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2392 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_22
timestamp 1679235063
transform 1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1679235063
transform 1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_35
timestamp 1679235063
transform 1 0 4324 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1679235063
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_59
timestamp 1679235063
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_70
timestamp 1679235063
transform 1 0 7544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1679235063
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1679235063
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1679235063
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_163
timestamp 1679235063
transform 1 0 16100 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1679235063
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_179
timestamp 1679235063
transform 1 0 17572 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_186
timestamp 1679235063
transform 1 0 18216 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1679235063
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1679235063
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1679235063
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1679235063
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_15
timestamp 1679235063
transform 1 0 2484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1679235063
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_77
timestamp 1679235063
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_81
timestamp 1679235063
transform 1 0 8556 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1679235063
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_113
timestamp 1679235063
transform 1 0 11500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1679235063
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_122
timestamp 1679235063
transform 1 0 12328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_135
timestamp 1679235063
transform 1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1679235063
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1679235063
transform 1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_175
timestamp 1679235063
transform 1 0 17204 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_179
timestamp 1679235063
transform 1 0 17572 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_192
timestamp 1679235063
transform 1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_200
timestamp 1679235063
transform 1 0 19504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_213
timestamp 1679235063
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_220
timestamp 1679235063
transform 1 0 21344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_230
timestamp 1679235063
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1679235063
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_15
timestamp 1679235063
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1679235063
transform 1 0 3680 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_42
timestamp 1679235063
transform 1 0 4968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1679235063
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1679235063
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1679235063
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1679235063
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1679235063
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 1679235063
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1679235063
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1679235063
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_171
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_182
timestamp 1679235063
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_194
timestamp 1679235063
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1679235063
transform 1 0 19504 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1679235063
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1679235063
transform 1 0 22264 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_241
timestamp 1679235063
transform 1 0 23276 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_245
timestamp 1679235063
transform 1 0 23644 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1679235063
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1679235063
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_47
timestamp 1679235063
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_54
timestamp 1679235063
transform 1 0 6072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1679235063
transform 1 0 6624 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_70
timestamp 1679235063
transform 1 0 7544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_96
timestamp 1679235063
transform 1 0 9936 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_100
timestamp 1679235063
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_125
timestamp 1679235063
transform 1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1679235063
transform 1 0 14444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_155
timestamp 1679235063
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_160
timestamp 1679235063
transform 1 0 15824 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_166
timestamp 1679235063
transform 1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1679235063
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_183
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1679235063
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_203
timestamp 1679235063
transform 1 0 19780 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_208
timestamp 1679235063
transform 1 0 20240 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1679235063
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1679235063
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1679235063
transform 1 0 3588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_32
timestamp 1679235063
transform 1 0 4048 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_40
timestamp 1679235063
transform 1 0 4784 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1679235063
transform 1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1679235063
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1679235063
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1679235063
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_127
timestamp 1679235063
transform 1 0 12788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_137
timestamp 1679235063
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_141
timestamp 1679235063
transform 1 0 14076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1679235063
transform 1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1679235063
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1679235063
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_203
timestamp 1679235063
transform 1 0 19780 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_210
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_235
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_240
timestamp 1679235063
transform 1 0 23184 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1679235063
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1679235063
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_35
timestamp 1679235063
transform 1 0 4324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1679235063
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_54
timestamp 1679235063
transform 1 0 6072 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1679235063
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1679235063
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_101
timestamp 1679235063
transform 1 0 10396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_114
timestamp 1679235063
transform 1 0 11592 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1679235063
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1679235063
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1679235063
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1679235063
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_187
timestamp 1679235063
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1679235063
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_216
timestamp 1679235063
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_220
timestamp 1679235063
transform 1 0 21344 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1679235063
transform 1 0 21712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1679235063
transform 1 0 22080 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1679235063
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1679235063
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1679235063
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_44
timestamp 1679235063
transform 1 0 5152 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_63
timestamp 1679235063
transform 1 0 6900 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1679235063
transform 1 0 9200 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1679235063
transform 1 0 10396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_105
timestamp 1679235063
transform 1 0 10764 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_119
timestamp 1679235063
transform 1 0 12052 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_130
timestamp 1679235063
transform 1 0 13064 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1679235063
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_161
timestamp 1679235063
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1679235063
transform 1 0 17572 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1679235063
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1679235063
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_247
timestamp 1679235063
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_260
timestamp 1679235063
transform 1 0 25024 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1679235063
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_45
timestamp 1679235063
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1679235063
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_69
timestamp 1679235063
transform 1 0 7452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1679235063
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_117
timestamp 1679235063
transform 1 0 11868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_121
timestamp 1679235063
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_133
timestamp 1679235063
transform 1 0 13340 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_137
timestamp 1679235063
transform 1 0 13708 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1679235063
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_162
timestamp 1679235063
transform 1 0 16008 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1679235063
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_178
timestamp 1679235063
transform 1 0 17480 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_188
timestamp 1679235063
transform 1 0 18400 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1679235063
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1679235063
transform 1 0 20516 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1679235063
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_263
timestamp 1679235063
transform 1 0 25300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_27
timestamp 1679235063
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1679235063
transform 1 0 4140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_42
timestamp 1679235063
transform 1 0 4968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1679235063
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_70
timestamp 1679235063
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_76
timestamp 1679235063
transform 1 0 8096 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_100
timestamp 1679235063
transform 1 0 10304 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_104
timestamp 1679235063
transform 1 0 10672 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1679235063
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1679235063
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1679235063
transform 1 0 14168 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_192
timestamp 1679235063
transform 1 0 18768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_199
timestamp 1679235063
transform 1 0 19412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1679235063
transform 1 0 20424 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1679235063
transform 1 0 22816 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_242
timestamp 1679235063
transform 1 0 23368 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1679235063
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_41
timestamp 1679235063
transform 1 0 4876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_44
timestamp 1679235063
transform 1 0 5152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1679235063
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1679235063
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1679235063
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1679235063
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1679235063
transform 1 0 14444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1679235063
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_167
timestamp 1679235063
transform 1 0 16468 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_179
timestamp 1679235063
transform 1 0 17572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_191
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1679235063
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1679235063
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1679235063
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_228
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_232
timestamp 1679235063
transform 1 0 22448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1679235063
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1679235063
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1679235063
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1679235063
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_43
timestamp 1679235063
transform 1 0 5060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_59
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_70
timestamp 1679235063
transform 1 0 7544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_82
timestamp 1679235063
transform 1 0 8648 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_88
timestamp 1679235063
transform 1 0 9200 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1679235063
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_124
timestamp 1679235063
transform 1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_148
timestamp 1679235063
transform 1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_160
timestamp 1679235063
transform 1 0 15824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1679235063
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_199
timestamp 1679235063
transform 1 0 19412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_204
timestamp 1679235063
transform 1 0 19872 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_260
timestamp 1679235063
transform 1 0 25024 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1679235063
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1679235063
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1679235063
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1679235063
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1679235063
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1679235063
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_112
timestamp 1679235063
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_115
timestamp 1679235063
transform 1 0 11684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1679235063
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_147
timestamp 1679235063
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1679235063
transform 1 0 15548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_170
timestamp 1679235063
transform 1 0 16744 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_182
timestamp 1679235063
transform 1 0 17848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_201
timestamp 1679235063
transform 1 0 19596 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_212
timestamp 1679235063
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1679235063
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_241
timestamp 1679235063
transform 1 0 23276 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_245
timestamp 1679235063
transform 1 0 23644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1679235063
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1679235063
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1679235063
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1679235063
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1679235063
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1679235063
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_63
timestamp 1679235063
transform 1 0 6900 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1679235063
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1679235063
transform 1 0 10396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_105
timestamp 1679235063
transform 1 0 10764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1679235063
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1679235063
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_160
timestamp 1679235063
transform 1 0 15824 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1679235063
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_192
timestamp 1679235063
transform 1 0 18768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_198
timestamp 1679235063
transform 1 0 19320 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_209
timestamp 1679235063
transform 1 0 20332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1679235063
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1679235063
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1679235063
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1679235063
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1679235063
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_63
timestamp 1679235063
transform 1 0 6900 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_70
timestamp 1679235063
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_107
timestamp 1679235063
transform 1 0 10948 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_124
timestamp 1679235063
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1679235063
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1679235063
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_176
timestamp 1679235063
transform 1 0 17296 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_184
timestamp 1679235063
transform 1 0 18032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_201
timestamp 1679235063
transform 1 0 19596 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_213
timestamp 1679235063
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_225
timestamp 1679235063
transform 1 0 21804 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_231
timestamp 1679235063
transform 1 0 22356 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1679235063
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1679235063
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1679235063
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1679235063
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1679235063
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_60
timestamp 1679235063
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_73
timestamp 1679235063
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_79
timestamp 1679235063
transform 1 0 8372 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_96
timestamp 1679235063
transform 1 0 9936 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_119
timestamp 1679235063
transform 1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1679235063
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_144
timestamp 1679235063
transform 1 0 14352 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_156
timestamp 1679235063
transform 1 0 15456 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1679235063
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1679235063
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1679235063
transform 1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1679235063
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_215
timestamp 1679235063
transform 1 0 20884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1679235063
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1679235063
transform 1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1679235063
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1679235063
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1679235063
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 1679235063
transform 1 0 5612 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_58
timestamp 1679235063
transform 1 0 6440 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1679235063
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1679235063
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_93
timestamp 1679235063
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1679235063
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1679235063
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1679235063
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_151
timestamp 1679235063
transform 1 0 14996 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_159
timestamp 1679235063
transform 1 0 15732 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1679235063
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_208
timestamp 1679235063
transform 1 0 20240 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_212
timestamp 1679235063
transform 1 0 20608 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_223
timestamp 1679235063
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_247
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1679235063
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_263
timestamp 1679235063
transform 1 0 25300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1679235063
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1679235063
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1679235063
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1679235063
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1679235063
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_77
timestamp 1679235063
transform 1 0 8188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_101
timestamp 1679235063
transform 1 0 10396 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1679235063
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1679235063
transform 1 0 12420 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_136
timestamp 1679235063
transform 1 0 13616 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_149
timestamp 1679235063
transform 1 0 14812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_161
timestamp 1679235063
transform 1 0 15916 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_165
timestamp 1679235063
transform 1 0 16284 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_180
timestamp 1679235063
transform 1 0 17664 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_186
timestamp 1679235063
transform 1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_198
timestamp 1679235063
transform 1 0 19320 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1679235063
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_229
timestamp 1679235063
transform 1 0 22172 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_240
timestamp 1679235063
transform 1 0 23184 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1679235063
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1679235063
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1679235063
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1679235063
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1679235063
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_65
timestamp 1679235063
transform 1 0 7084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_73
timestamp 1679235063
transform 1 0 7820 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1679235063
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1679235063
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_131
timestamp 1679235063
transform 1 0 13156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1679235063
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_154
timestamp 1679235063
transform 1 0 15272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_167
timestamp 1679235063
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_171
timestamp 1679235063
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1679235063
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_192
timestamp 1679235063
transform 1 0 18768 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_197
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1679235063
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_216
timestamp 1679235063
transform 1 0 20976 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_220
timestamp 1679235063
transform 1 0 21344 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1679235063
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1679235063
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_263
timestamp 1679235063
transform 1 0 25300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1679235063
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1679235063
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1679235063
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1679235063
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1679235063
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_65
timestamp 1679235063
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_74
timestamp 1679235063
transform 1 0 7912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_86
timestamp 1679235063
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1679235063
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_123
timestamp 1679235063
transform 1 0 12420 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_147
timestamp 1679235063
transform 1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_160
timestamp 1679235063
transform 1 0 15824 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1679235063
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_193
timestamp 1679235063
transform 1 0 18860 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_197
timestamp 1679235063
transform 1 0 19228 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_208
timestamp 1679235063
transform 1 0 20240 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_220
timestamp 1679235063
transform 1 0 21344 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1679235063
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1679235063
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_259
timestamp 1679235063
transform 1 0 24932 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_263
timestamp 1679235063
transform 1 0 25300 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1679235063
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1679235063
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1679235063
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_53
timestamp 1679235063
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_61
timestamp 1679235063
transform 1 0 6716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_70
timestamp 1679235063
transform 1 0 7544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1679235063
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_91
timestamp 1679235063
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_103
timestamp 1679235063
transform 1 0 10580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_115
timestamp 1679235063
transform 1 0 11684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_128
timestamp 1679235063
transform 1 0 12880 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_134
timestamp 1679235063
transform 1 0 13432 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1679235063
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_143
timestamp 1679235063
transform 1 0 14260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_154
timestamp 1679235063
transform 1 0 15272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp 1679235063
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_178
timestamp 1679235063
transform 1 0 17480 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_182
timestamp 1679235063
transform 1 0 17848 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_191
timestamp 1679235063
transform 1 0 18676 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1679235063
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_219
timestamp 1679235063
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_226
timestamp 1679235063
transform 1 0 21896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1679235063
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1679235063
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1679235063
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1679235063
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1679235063
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1679235063
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1679235063
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1679235063
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_77
timestamp 1679235063
transform 1 0 8188 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1679235063
transform 1 0 9016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1679235063
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1679235063
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1679235063
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_138
timestamp 1679235063
transform 1 0 13800 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_146
timestamp 1679235063
transform 1 0 14536 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_157
timestamp 1679235063
transform 1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_161
timestamp 1679235063
transform 1 0 15916 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1679235063
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_179
timestamp 1679235063
transform 1 0 17572 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_183
timestamp 1679235063
transform 1 0 17940 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_204
timestamp 1679235063
transform 1 0 19872 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_216
timestamp 1679235063
transform 1 0 20976 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_220
timestamp 1679235063
transform 1 0 21344 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_247
timestamp 1679235063
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_253
timestamp 1679235063
transform 1 0 24380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_263
timestamp 1679235063
transform 1 0 25300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1679235063
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1679235063
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1679235063
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1679235063
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1679235063
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1679235063
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1679235063
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_88
timestamp 1679235063
transform 1 0 9200 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_94
timestamp 1679235063
transform 1 0 9752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_115
timestamp 1679235063
transform 1 0 11684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_121
timestamp 1679235063
transform 1 0 12236 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_126
timestamp 1679235063
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1679235063
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_147
timestamp 1679235063
transform 1 0 14628 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_158
timestamp 1679235063
transform 1 0 15640 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_171
timestamp 1679235063
transform 1 0 16836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_184
timestamp 1679235063
transform 1 0 18032 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1679235063
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_207
timestamp 1679235063
transform 1 0 20148 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_211
timestamp 1679235063
transform 1 0 20516 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_232
timestamp 1679235063
transform 1 0 22448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_245
timestamp 1679235063
transform 1 0 23644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_249
timestamp 1679235063
transform 1 0 24012 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp 1679235063
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1679235063
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1679235063
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1679235063
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1679235063
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1679235063
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1679235063
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_81
timestamp 1679235063
transform 1 0 8556 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_102
timestamp 1679235063
transform 1 0 10488 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_106
timestamp 1679235063
transform 1 0 10856 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_136
timestamp 1679235063
transform 1 0 13616 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_160
timestamp 1679235063
transform 1 0 15824 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_164
timestamp 1679235063
transform 1 0 16192 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1679235063
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_175
timestamp 1679235063
transform 1 0 17204 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_199
timestamp 1679235063
transform 1 0 19412 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_211
timestamp 1679235063
transform 1 0 20516 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_215
timestamp 1679235063
transform 1 0 20884 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1679235063
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_247
timestamp 1679235063
transform 1 0 23828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_252
timestamp 1679235063
transform 1 0 24288 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_264
timestamp 1679235063
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1679235063
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1679235063
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1679235063
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_65
timestamp 1679235063
transform 1 0 7084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_73
timestamp 1679235063
transform 1 0 7820 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1679235063
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_102
timestamp 1679235063
transform 1 0 10488 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_128
timestamp 1679235063
transform 1 0 12880 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_132
timestamp 1679235063
transform 1 0 13248 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1679235063
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_152
timestamp 1679235063
transform 1 0 15088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_165
timestamp 1679235063
transform 1 0 16284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_178
timestamp 1679235063
transform 1 0 17480 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_191
timestamp 1679235063
transform 1 0 18676 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1679235063
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1679235063
transform 1 0 20424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_225
timestamp 1679235063
transform 1 0 21804 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_238
timestamp 1679235063
transform 1 0 23000 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_248
timestamp 1679235063
transform 1 0 23920 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1679235063
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1679235063
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1679235063
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1679235063
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1679235063
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1679235063
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1679235063
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1679235063
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1679235063
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_89
timestamp 1679235063
transform 1 0 9292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1679235063
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_116
timestamp 1679235063
transform 1 0 11776 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_126
timestamp 1679235063
transform 1 0 12696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_150
timestamp 1679235063
transform 1 0 14904 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_154
timestamp 1679235063
transform 1 0 15272 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1679235063
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1679235063
transform 1 0 17572 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_191
timestamp 1679235063
transform 1 0 18676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_199
timestamp 1679235063
transform 1 0 19412 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_210
timestamp 1679235063
transform 1 0 20424 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1679235063
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_236
timestamp 1679235063
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_249
timestamp 1679235063
transform 1 0 24012 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_261
timestamp 1679235063
transform 1 0 25116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_265
timestamp 1679235063
transform 1 0 25484 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1679235063
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1679235063
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1679235063
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1679235063
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1679235063
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1679235063
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_97
timestamp 1679235063
transform 1 0 10028 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_106
timestamp 1679235063
transform 1 0 10856 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_130
timestamp 1679235063
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_134
timestamp 1679235063
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1679235063
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_141
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_147
timestamp 1679235063
transform 1 0 14628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_160
timestamp 1679235063
transform 1 0 15824 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_164
timestamp 1679235063
transform 1 0 16192 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1679235063
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1679235063
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1679235063
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1679235063
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_225
timestamp 1679235063
transform 1 0 21804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_237
timestamp 1679235063
transform 1 0 22908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1679235063
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_263
timestamp 1679235063
transform 1 0 25300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1679235063
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1679235063
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1679235063
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1679235063
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1679235063
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_85
timestamp 1679235063
transform 1 0 8924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_94
timestamp 1679235063
transform 1 0 9752 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1679235063
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_145
timestamp 1679235063
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_160
timestamp 1679235063
transform 1 0 15824 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_180
timestamp 1679235063
transform 1 0 17664 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_192
timestamp 1679235063
transform 1 0 18768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1679235063
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 1679235063
transform 1 0 19780 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_213
timestamp 1679235063
transform 1 0 20700 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1679235063
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_231
timestamp 1679235063
transform 1 0 22356 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_255
timestamp 1679235063
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1679235063
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1679235063
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1679235063
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1679235063
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1679235063
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1679235063
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1679235063
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1679235063
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_97
timestamp 1679235063
transform 1 0 10028 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_111
timestamp 1679235063
transform 1 0 11316 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_123
timestamp 1679235063
transform 1 0 12420 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_135
timestamp 1679235063
transform 1 0 13524 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_154
timestamp 1679235063
transform 1 0 15272 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_158
timestamp 1679235063
transform 1 0 15640 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1679235063
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1679235063
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_207
timestamp 1679235063
transform 1 0 20148 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_213
timestamp 1679235063
transform 1 0 20700 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_237
timestamp 1679235063
transform 1 0 22908 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1679235063
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_263
timestamp 1679235063
transform 1 0 25300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1679235063
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1679235063
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1679235063
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1679235063
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1679235063
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1679235063
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1679235063
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_93
timestamp 1679235063
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_101
timestamp 1679235063
transform 1 0 10396 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1679235063
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_129
timestamp 1679235063
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_141
timestamp 1679235063
transform 1 0 14076 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_145
timestamp 1679235063
transform 1 0 14444 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1679235063
transform 1 0 15272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1679235063
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_174
timestamp 1679235063
transform 1 0 17112 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_184
timestamp 1679235063
transform 1 0 18032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1679235063
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_200
timestamp 1679235063
transform 1 0 19504 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_204
timestamp 1679235063
transform 1 0 19872 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_217
timestamp 1679235063
transform 1 0 21068 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_221
timestamp 1679235063
transform 1 0 21436 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_235
timestamp 1679235063
transform 1 0 22724 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_241
timestamp 1679235063
transform 1 0 23276 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_262
timestamp 1679235063
transform 1 0 25208 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1679235063
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1679235063
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1679235063
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1679235063
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1679235063
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_96
timestamp 1679235063
transform 1 0 9936 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_108
timestamp 1679235063
transform 1 0 11040 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_114
timestamp 1679235063
transform 1 0 11592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_123
timestamp 1679235063
transform 1 0 12420 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_127
timestamp 1679235063
transform 1 0 12788 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1679235063
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_163
timestamp 1679235063
transform 1 0 16100 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_168
timestamp 1679235063
transform 1 0 16560 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_171
timestamp 1679235063
transform 1 0 16836 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 1679235063
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_219
timestamp 1679235063
transform 1 0 21252 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_225
timestamp 1679235063
transform 1 0 21804 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_236
timestamp 1679235063
transform 1 0 22816 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1679235063
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_263
timestamp 1679235063
transform 1 0 25300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1679235063
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1679235063
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1679235063
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1679235063
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1679235063
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1679235063
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1679235063
transform 1 0 8556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_85
timestamp 1679235063
transform 1 0 8924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_89
timestamp 1679235063
transform 1 0 9292 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_101
timestamp 1679235063
transform 1 0 10396 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 1679235063
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1679235063
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1679235063
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1679235063
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1679235063
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_173
timestamp 1679235063
transform 1 0 17020 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_179
timestamp 1679235063
transform 1 0 17572 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_200
timestamp 1679235063
transform 1 0 19504 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_215
timestamp 1679235063
transform 1 0 20884 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1679235063
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_238
timestamp 1679235063
transform 1 0 23000 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_262
timestamp 1679235063
transform 1 0 25208 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1679235063
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1679235063
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1679235063
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1679235063
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1679235063
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1679235063
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1679235063
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_92
timestamp 1679235063
transform 1 0 9568 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_104
timestamp 1679235063
transform 1 0 10672 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_116
timestamp 1679235063
transform 1 0 11776 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_128
timestamp 1679235063
transform 1 0 12880 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_153
timestamp 1679235063
transform 1 0 15180 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_164
timestamp 1679235063
transform 1 0 16192 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_177
timestamp 1679235063
transform 1 0 17388 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_189
timestamp 1679235063
transform 1 0 18492 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1679235063
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_219
timestamp 1679235063
transform 1 0 21252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_226
timestamp 1679235063
transform 1 0 21896 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1679235063
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1679235063
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1679235063
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1679235063
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1679235063
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1679235063
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1679235063
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1679235063
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1679235063
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1679235063
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1679235063
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1679235063
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1679235063
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1679235063
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1679235063
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1679235063
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_161
timestamp 1679235063
transform 1 0 15916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_177
timestamp 1679235063
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_186
timestamp 1679235063
transform 1 0 18216 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_191
timestamp 1679235063
transform 1 0 18676 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_196
timestamp 1679235063
transform 1 0 19136 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_220
timestamp 1679235063
transform 1 0 21344 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1679235063
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_260
timestamp 1679235063
transform 1 0 25024 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1679235063
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1679235063
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1679235063
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1679235063
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1679235063
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1679235063
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1679235063
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_93
timestamp 1679235063
transform 1 0 9660 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1679235063
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1679235063
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1679235063
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1679235063
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_141
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_155
timestamp 1679235063
transform 1 0 15364 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_159
timestamp 1679235063
transform 1 0 15732 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_171
timestamp 1679235063
transform 1 0 16836 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_181
timestamp 1679235063
transform 1 0 17756 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1679235063
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1679235063
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_243
timestamp 1679235063
transform 1 0 23460 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1679235063
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_263
timestamp 1679235063
transform 1 0 25300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1679235063
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1679235063
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1679235063
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1679235063
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1679235063
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1679235063
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1679235063
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1679235063
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1679235063
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1679235063
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1679235063
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1679235063
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1679235063
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_181
timestamp 1679235063
transform 1 0 17756 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_185
timestamp 1679235063
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_197
timestamp 1679235063
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1679235063
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1679235063
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1679235063
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_247
timestamp 1679235063
transform 1 0 23828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_259
timestamp 1679235063
transform 1 0 24932 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_265
timestamp 1679235063
transform 1 0 25484 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1679235063
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1679235063
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1679235063
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1679235063
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1679235063
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1679235063
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1679235063
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1679235063
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1679235063
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1679235063
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1679235063
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1679235063
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_177
timestamp 1679235063
transform 1 0 17388 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_187
timestamp 1679235063
transform 1 0 18308 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1679235063
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_199
timestamp 1679235063
transform 1 0 19412 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_209
timestamp 1679235063
transform 1 0 20332 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_221
timestamp 1679235063
transform 1 0 21436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_226
timestamp 1679235063
transform 1 0 21896 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1679235063
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_244
timestamp 1679235063
transform 1 0 23552 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_263
timestamp 1679235063
transform 1 0 25300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1679235063
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1679235063
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1679235063
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1679235063
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1679235063
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1679235063
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_81
timestamp 1679235063
transform 1 0 8556 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_86
timestamp 1679235063
transform 1 0 9016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1679235063
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_117
timestamp 1679235063
transform 1 0 11868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_129
timestamp 1679235063
transform 1 0 12972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1679235063
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1679235063
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1679235063
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1679235063
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_193
timestamp 1679235063
transform 1 0 18860 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_209
timestamp 1679235063
transform 1 0 20332 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1679235063
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1679235063
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1679235063
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_260
timestamp 1679235063
transform 1 0 25024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1679235063
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1679235063
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1679235063
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1679235063
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1679235063
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1679235063
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1679235063
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1679235063
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1679235063
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1679235063
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1679235063
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1679235063
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1679235063
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1679235063
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1679235063
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1679235063
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_213
timestamp 1679235063
transform 1 0 20700 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_225
timestamp 1679235063
transform 1 0 21804 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1679235063
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1679235063
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_263
timestamp 1679235063
transform 1 0 25300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1679235063
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1679235063
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1679235063
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1679235063
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1679235063
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1679235063
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1679235063
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1679235063
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1679235063
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1679235063
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1679235063
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1679235063
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1679235063
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1679235063
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1679235063
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_205
timestamp 1679235063
transform 1 0 19964 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_213
timestamp 1679235063
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1679235063
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_229
timestamp 1679235063
transform 1 0 22172 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_238
timestamp 1679235063
transform 1 0 23000 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_252
timestamp 1679235063
transform 1 0 24288 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1679235063
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1679235063
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1679235063
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1679235063
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1679235063
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1679235063
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1679235063
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1679235063
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1679235063
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1679235063
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1679235063
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1679235063
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1679235063
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1679235063
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1679235063
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1679235063
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1679235063
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_221
timestamp 1679235063
transform 1 0 21436 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_229
timestamp 1679235063
transform 1 0 22172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1679235063
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1679235063
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_263
timestamp 1679235063
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1679235063
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1679235063
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1679235063
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1679235063
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1679235063
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1679235063
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1679235063
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1679235063
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1679235063
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1679235063
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1679235063
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1679235063
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1679235063
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_123
timestamp 1679235063
transform 1 0 12420 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_135
timestamp 1679235063
transform 1 0 13524 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_147
timestamp 1679235063
transform 1 0 14628 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_159
timestamp 1679235063
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1679235063
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1679235063
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1679235063
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1679235063
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1679235063
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1679235063
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1679235063
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_225
timestamp 1679235063
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_233
timestamp 1679235063
transform 1 0 22540 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_245
timestamp 1679235063
transform 1 0 23644 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_257
timestamp 1679235063
transform 1 0 24748 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_261
timestamp 1679235063
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_265
timestamp 1679235063
transform 1 0 25484 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1679235063
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1679235063
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1679235063
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1679235063
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1679235063
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1679235063
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1679235063
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1679235063
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1679235063
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1679235063
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1679235063
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1679235063
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1679235063
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1679235063
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1679235063
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1679235063
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1679235063
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1679235063
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_177
timestamp 1679235063
transform 1 0 17388 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_185
timestamp 1679235063
transform 1 0 18124 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1679235063
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1679235063
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1679235063
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1679235063
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_233
timestamp 1679235063
transform 1 0 22540 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_241
timestamp 1679235063
transform 1 0 23276 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_245
timestamp 1679235063
transform 1 0 23644 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1679235063
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1679235063
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_263
timestamp 1679235063
transform 1 0 25300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1679235063
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1679235063
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1679235063
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1679235063
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1679235063
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1679235063
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1679235063
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1679235063
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_84
timestamp 1679235063
transform 1 0 8832 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_96
timestamp 1679235063
transform 1 0 9936 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_108
timestamp 1679235063
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1679235063
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1679235063
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1679235063
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1679235063
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1679235063
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1679235063
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1679235063
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1679235063
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1679235063
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1679235063
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1679235063
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1679235063
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1679235063
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1679235063
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_252
timestamp 1679235063
transform 1 0 24288 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_264
timestamp 1679235063
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1679235063
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1679235063
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1679235063
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1679235063
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1679235063
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1679235063
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1679235063
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1679235063
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1679235063
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1679235063
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1679235063
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_109
timestamp 1679235063
transform 1 0 11132 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_118
timestamp 1679235063
transform 1 0 11960 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_130
timestamp 1679235063
transform 1 0 13064 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_138
timestamp 1679235063
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1679235063
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1679235063
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1679235063
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1679235063
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1679235063
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1679235063
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1679235063
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1679235063
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1679235063
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1679235063
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_245
timestamp 1679235063
transform 1 0 23644 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_249
timestamp 1679235063
transform 1 0 24012 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_255
timestamp 1679235063
transform 1 0 24564 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_258
timestamp 1679235063
transform 1 0 24840 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1679235063
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1679235063
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1679235063
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1679235063
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1679235063
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1679235063
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1679235063
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1679235063
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1679235063
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1679235063
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1679235063
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1679235063
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1679235063
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1679235063
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1679235063
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1679235063
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1679235063
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1679235063
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1679235063
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1679235063
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1679235063
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1679235063
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1679235063
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1679235063
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1679235063
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1679235063
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1679235063
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_249
timestamp 1679235063
transform 1 0 24012 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_256
timestamp 1679235063
transform 1 0 24656 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1679235063
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1679235063
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1679235063
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1679235063
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1679235063
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1679235063
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1679235063
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1679235063
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1679235063
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1679235063
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1679235063
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1679235063
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1679235063
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1679235063
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1679235063
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1679235063
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1679235063
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1679235063
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1679235063
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1679235063
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1679235063
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1679235063
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1679235063
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1679235063
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1679235063
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1679235063
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1679235063
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1679235063
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1679235063
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_259
timestamp 1679235063
transform 1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_264
timestamp 1679235063
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1679235063
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1679235063
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1679235063
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1679235063
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1679235063
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1679235063
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1679235063
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1679235063
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1679235063
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1679235063
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1679235063
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1679235063
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1679235063
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1679235063
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1679235063
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1679235063
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1679235063
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1679235063
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1679235063
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1679235063
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_193
timestamp 1679235063
transform 1 0 18860 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_207
timestamp 1679235063
transform 1 0 20148 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_219
timestamp 1679235063
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1679235063
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1679235063
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1679235063
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_249
timestamp 1679235063
transform 1 0 24012 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_252
timestamp 1679235063
transform 1 0 24288 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_257
timestamp 1679235063
transform 1 0 24748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1679235063
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1679235063
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1679235063
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1679235063
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1679235063
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1679235063
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1679235063
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1679235063
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1679235063
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1679235063
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1679235063
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1679235063
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1679235063
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1679235063
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1679235063
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1679235063
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1679235063
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1679235063
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1679235063
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1679235063
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1679235063
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1679235063
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1679235063
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1679235063
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1679235063
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1679235063
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1679235063
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1679235063
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_253
timestamp 1679235063
transform 1 0 24380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_258
timestamp 1679235063
transform 1 0 24840 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1679235063
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1679235063
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1679235063
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1679235063
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1679235063
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1679235063
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1679235063
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1679235063
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1679235063
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1679235063
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1679235063
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1679235063
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1679235063
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1679235063
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1679235063
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1679235063
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1679235063
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1679235063
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1679235063
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1679235063
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1679235063
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1679235063
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1679235063
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1679235063
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1679235063
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1679235063
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1679235063
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1679235063
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_261
timestamp 1679235063
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1679235063
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1679235063
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1679235063
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1679235063
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1679235063
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1679235063
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1679235063
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1679235063
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1679235063
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1679235063
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_113
timestamp 1679235063
transform 1 0 11500 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_119
timestamp 1679235063
transform 1 0 12052 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_131
timestamp 1679235063
transform 1 0 13156 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1679235063
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1679235063
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1679235063
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1679235063
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1679235063
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1679235063
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1679235063
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1679235063
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1679235063
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1679235063
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1679235063
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1679235063
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1679235063
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1679235063
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1679235063
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1679235063
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1679235063
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1679235063
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1679235063
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1679235063
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1679235063
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1679235063
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1679235063
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1679235063
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1679235063
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1679235063
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1679235063
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1679235063
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1679235063
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1679235063
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1679235063
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1679235063
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1679235063
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1679235063
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1679235063
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1679235063
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1679235063
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1679235063
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1679235063
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1679235063
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1679235063
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1679235063
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1679235063
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_257
timestamp 1679235063
transform 1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1679235063
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1679235063
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1679235063
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1679235063
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1679235063
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1679235063
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1679235063
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1679235063
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1679235063
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1679235063
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1679235063
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_93
timestamp 1679235063
transform 1 0 9660 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_104
timestamp 1679235063
transform 1 0 10672 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_116
timestamp 1679235063
transform 1 0 11776 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_128
timestamp 1679235063
transform 1 0 12880 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1679235063
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1679235063
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1679235063
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1679235063
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1679235063
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1679235063
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1679235063
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_209
timestamp 1679235063
transform 1 0 20332 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_231
timestamp 1679235063
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_235
timestamp 1679235063
transform 1 0 22724 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_247
timestamp 1679235063
transform 1 0 23828 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1679235063
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1679235063
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_261
timestamp 1679235063
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1679235063
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1679235063
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1679235063
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1679235063
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1679235063
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1679235063
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1679235063
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1679235063
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1679235063
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_93
timestamp 1679235063
transform 1 0 9660 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_107
timestamp 1679235063
transform 1 0 10948 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1679235063
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_115
timestamp 1679235063
transform 1 0 11684 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_127
timestamp 1679235063
transform 1 0 12788 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_139
timestamp 1679235063
transform 1 0 13892 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_151
timestamp 1679235063
transform 1 0 14996 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_163
timestamp 1679235063
transform 1 0 16100 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1679235063
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1679235063
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1679235063
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1679235063
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1679235063
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1679235063
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1679235063
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1679235063
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1679235063
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_249
timestamp 1679235063
transform 1 0 24012 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_255
timestamp 1679235063
transform 1 0 24564 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_258
timestamp 1679235063
transform 1 0 24840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1679235063
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1679235063
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1679235063
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1679235063
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1679235063
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1679235063
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1679235063
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1679235063
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1679235063
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1679235063
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1679235063
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_107
timestamp 1679235063
transform 1 0 10948 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_119
timestamp 1679235063
transform 1 0 12052 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_131
timestamp 1679235063
transform 1 0 13156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1679235063
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1679235063
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1679235063
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1679235063
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1679235063
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1679235063
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1679235063
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1679235063
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1679235063
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1679235063
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1679235063
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1679235063
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1679235063
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1679235063
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1679235063
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1679235063
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1679235063
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1679235063
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1679235063
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1679235063
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1679235063
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1679235063
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1679235063
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_81
timestamp 1679235063
transform 1 0 8556 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_110
timestamp 1679235063
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1679235063
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_122
timestamp 1679235063
transform 1 0 12328 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_126
timestamp 1679235063
transform 1 0 12696 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_138
timestamp 1679235063
transform 1 0 13800 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_150
timestamp 1679235063
transform 1 0 14904 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_162
timestamp 1679235063
transform 1 0 16008 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1679235063
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1679235063
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1679235063
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1679235063
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1679235063
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1679235063
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1679235063
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1679235063
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1679235063
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_261
timestamp 1679235063
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1679235063
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1679235063
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1679235063
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1679235063
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1679235063
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1679235063
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1679235063
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1679235063
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1679235063
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1679235063
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_95
timestamp 1679235063
transform 1 0 9844 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_124
timestamp 1679235063
transform 1 0 12512 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1679235063
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1679235063
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_153
timestamp 1679235063
transform 1 0 15180 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_178
timestamp 1679235063
transform 1 0 17480 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_190
timestamp 1679235063
transform 1 0 18584 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1679235063
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1679235063
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1679235063
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1679235063
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1679235063
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1679235063
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1679235063
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_259
timestamp 1679235063
transform 1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1679235063
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1679235063
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1679235063
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1679235063
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1679235063
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1679235063
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1679235063
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1679235063
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1679235063
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1679235063
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1679235063
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1679235063
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1679235063
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_113
timestamp 1679235063
transform 1 0 11500 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_119
timestamp 1679235063
transform 1 0 12052 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_141
timestamp 1679235063
transform 1 0 14076 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1679235063
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1679235063
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1679235063
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1679235063
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1679235063
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1679235063
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1679235063
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1679235063
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1679235063
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1679235063
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1679235063
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1679235063
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1679235063
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1679235063
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1679235063
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1679235063
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1679235063
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1679235063
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1679235063
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1679235063
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1679235063
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_95
timestamp 1679235063
transform 1 0 9844 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_106
timestamp 1679235063
transform 1 0 10856 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_110
timestamp 1679235063
transform 1 0 11224 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_122
timestamp 1679235063
transform 1 0 12328 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_130
timestamp 1679235063
transform 1 0 13064 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1679235063
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1679235063
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1679235063
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_164
timestamp 1679235063
transform 1 0 16192 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_176
timestamp 1679235063
transform 1 0 17296 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_188
timestamp 1679235063
transform 1 0 18400 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1679235063
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1679235063
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1679235063
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_233
timestamp 1679235063
transform 1 0 22540 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_242
timestamp 1679235063
transform 1 0 23368 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1679235063
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1679235063
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1679235063
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1679235063
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1679235063
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1679235063
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1679235063
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1679235063
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1679235063
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1679235063
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_69
timestamp 1679235063
transform 1 0 7452 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_77
timestamp 1679235063
transform 1 0 8188 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_80
timestamp 1679235063
transform 1 0 8464 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_103
timestamp 1679235063
transform 1 0 10580 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1679235063
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_113
timestamp 1679235063
transform 1 0 11500 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_121
timestamp 1679235063
transform 1 0 12236 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_126
timestamp 1679235063
transform 1 0 12696 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_138
timestamp 1679235063
transform 1 0 13800 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_150
timestamp 1679235063
transform 1 0 14904 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_162
timestamp 1679235063
transform 1 0 16008 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1679235063
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1679235063
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1679235063
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1679235063
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1679235063
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1679235063
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1679235063
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1679235063
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1679235063
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_259
timestamp 1679235063
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1679235063
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1679235063
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1679235063
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1679235063
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1679235063
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1679235063
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_53
timestamp 1679235063
transform 1 0 5980 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_84_79
timestamp 1679235063
transform 1 0 8372 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1679235063
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_85
timestamp 1679235063
transform 1 0 8924 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_95
timestamp 1679235063
transform 1 0 9844 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_102
timestamp 1679235063
transform 1 0 10488 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_110
timestamp 1679235063
transform 1 0 11224 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_115
timestamp 1679235063
transform 1 0 11684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_127
timestamp 1679235063
transform 1 0 12788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1679235063
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1679235063
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1679235063
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1679235063
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1679235063
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1679235063
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1679235063
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1679235063
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1679235063
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1679235063
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1679235063
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1679235063
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1679235063
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1679235063
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1679235063
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1679235063
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1679235063
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1679235063
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1679235063
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1679235063
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1679235063
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1679235063
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1679235063
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_69
timestamp 1679235063
transform 1 0 7452 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_93
timestamp 1679235063
transform 1 0 9660 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_104
timestamp 1679235063
transform 1 0 10672 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_108
timestamp 1679235063
transform 1 0 11040 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1679235063
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1679235063
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1679235063
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1679235063
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1679235063
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1679235063
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1679235063
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1679235063
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1679235063
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1679235063
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1679235063
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1679235063
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1679235063
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1679235063
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1679235063
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1679235063
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1679235063
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1679235063
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1679235063
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1679235063
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1679235063
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1679235063
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1679235063
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1679235063
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1679235063
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1679235063
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1679235063
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1679235063
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1679235063
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1679235063
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1679235063
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1679235063
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1679235063
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1679235063
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1679235063
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1679235063
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1679235063
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1679235063
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1679235063
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1679235063
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_241
timestamp 1679235063
transform 1 0 23276 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_249
timestamp 1679235063
transform 1 0 24012 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1679235063
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1679235063
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1679235063
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1679235063
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1679235063
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1679235063
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1679235063
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1679235063
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1679235063
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1679235063
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1679235063
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1679235063
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1679235063
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1679235063
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1679235063
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1679235063
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1679235063
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1679235063
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1679235063
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1679235063
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1679235063
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1679235063
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1679235063
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1679235063
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1679235063
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1679235063
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1679235063
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1679235063
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1679235063
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1679235063
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1679235063
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1679235063
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1679235063
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1679235063
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1679235063
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1679235063
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1679235063
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1679235063
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1679235063
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1679235063
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1679235063
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1679235063
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1679235063
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1679235063
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1679235063
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1679235063
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1679235063
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1679235063
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1679235063
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1679235063
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1679235063
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1679235063
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1679235063
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1679235063
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1679235063
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1679235063
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1679235063
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1679235063
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1679235063
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1679235063
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1679235063
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1679235063
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1679235063
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1679235063
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1679235063
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1679235063
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1679235063
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1679235063
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_76
timestamp 1679235063
transform 1 0 8096 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_80
timestamp 1679235063
transform 1 0 8464 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_92
timestamp 1679235063
transform 1 0 9568 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_104
timestamp 1679235063
transform 1 0 10672 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1679235063
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1679235063
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1679235063
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1679235063
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1679235063
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1679235063
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1679235063
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1679235063
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1679235063
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1679235063
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1679235063
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1679235063
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1679235063
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1679235063
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1679235063
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_253
timestamp 1679235063
transform 1 0 24380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_256
timestamp 1679235063
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1679235063
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1679235063
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1679235063
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1679235063
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1679235063
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1679235063
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1679235063
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1679235063
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1679235063
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1679235063
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1679235063
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1679235063
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1679235063
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1679235063
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1679235063
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1679235063
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1679235063
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1679235063
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1679235063
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1679235063
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1679235063
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1679235063
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1679235063
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1679235063
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1679235063
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1679235063
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_245
timestamp 1679235063
transform 1 0 23644 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_253
timestamp 1679235063
transform 1 0 24380 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1679235063
transform 1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1679235063
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1679235063
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1679235063
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1679235063
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1679235063
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1679235063
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1679235063
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1679235063
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1679235063
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_81
timestamp 1679235063
transform 1 0 8556 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_86
timestamp 1679235063
transform 1 0 9016 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_98
timestamp 1679235063
transform 1 0 10120 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_110
timestamp 1679235063
transform 1 0 11224 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1679235063
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1679235063
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1679235063
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1679235063
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1679235063
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1679235063
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1679235063
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1679235063
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1679235063
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1679235063
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1679235063
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1679235063
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1679235063
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_245
timestamp 1679235063
transform 1 0 23644 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_249
timestamp 1679235063
transform 1 0 24012 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_254
timestamp 1679235063
transform 1 0 24472 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1679235063
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1679235063
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1679235063
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1679235063
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1679235063
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1679235063
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1679235063
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1679235063
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_92_74
timestamp 1679235063
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1679235063
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1679235063
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1679235063
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1679235063
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1679235063
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1679235063
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1679235063
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1679235063
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1679235063
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1679235063
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1679235063
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1679235063
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1679235063
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1679235063
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1679235063
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1679235063
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_233
timestamp 1679235063
transform 1 0 22540 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_242
timestamp 1679235063
transform 1 0 23368 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_250
timestamp 1679235063
transform 1 0 24104 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_253
timestamp 1679235063
transform 1 0 24380 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1679235063
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1679235063
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1679235063
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1679235063
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_39
timestamp 1679235063
transform 1 0 4692 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1679235063
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1679235063
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1679235063
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_62
timestamp 1679235063
transform 1 0 6808 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_74
timestamp 1679235063
transform 1 0 7912 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_86
timestamp 1679235063
transform 1 0 9016 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_98
timestamp 1679235063
transform 1 0 10120 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1679235063
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1679235063
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1679235063
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1679235063
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1679235063
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1679235063
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1679235063
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1679235063
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1679235063
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1679235063
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1679235063
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1679235063
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1679235063
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_225
timestamp 1679235063
transform 1 0 21804 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_233
timestamp 1679235063
transform 1 0 22540 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_239
timestamp 1679235063
transform 1 0 23092 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_251
timestamp 1679235063
transform 1 0 24196 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_263
timestamp 1679235063
transform 1 0 25300 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1679235063
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1679235063
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1679235063
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1679235063
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1679235063
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_61
timestamp 1679235063
transform 1 0 6716 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_73
timestamp 1679235063
transform 1 0 7820 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_81
timestamp 1679235063
transform 1 0 8556 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1679235063
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1679235063
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1679235063
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1679235063
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1679235063
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1679235063
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1679235063
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1679235063
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1679235063
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1679235063
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1679235063
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1679235063
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1679235063
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1679235063
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_221
timestamp 1679235063
transform 1 0 21436 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_229
timestamp 1679235063
transform 1 0 22172 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_235
timestamp 1679235063
transform 1 0 22724 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_247
timestamp 1679235063
transform 1 0 23828 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1679235063
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_263
timestamp 1679235063
transform 1 0 25300 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1679235063
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1679235063
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1679235063
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_29
timestamp 1679235063
transform 1 0 3772 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_47
timestamp 1679235063
transform 1 0 5428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1679235063
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_57
timestamp 1679235063
transform 1 0 6348 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_76
timestamp 1679235063
transform 1 0 8096 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_85
timestamp 1679235063
transform 1 0 8924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_97
timestamp 1679235063
transform 1 0 10028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_109
timestamp 1679235063
transform 1 0 11132 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1679235063
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_125
timestamp 1679235063
transform 1 0 12604 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_133
timestamp 1679235063
transform 1 0 13340 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1679235063
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_143
timestamp 1679235063
transform 1 0 14260 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1679235063
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_153
timestamp 1679235063
transform 1 0 15180 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_157
timestamp 1679235063
transform 1 0 15548 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1679235063
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1679235063
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_174
timestamp 1679235063
transform 1 0 17112 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_178
timestamp 1679235063
transform 1 0 17480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_183
timestamp 1679235063
transform 1 0 17940 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_187
timestamp 1679235063
transform 1 0 18308 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_193
timestamp 1679235063
transform 1 0 18860 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1679235063
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_209
timestamp 1679235063
transform 1 0 20332 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_217
timestamp 1679235063
transform 1 0 21068 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1679235063
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_227
timestamp 1679235063
transform 1 0 21988 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_238
timestamp 1679235063
transform 1 0 23000 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1679235063
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_253
timestamp 1679235063
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_263
timestamp 1679235063
transform 1 0 25300 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 24564 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 22540 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 24564 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold7
timestamp 1679235063
transform 1 0 21068 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold8
timestamp 1679235063
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 17940 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 11960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 14444 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 21988 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 19596 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 17480 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold17
timestamp 1679235063
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 7912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 12420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold21
timestamp 1679235063
transform 1 0 7268 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold22
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 9292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 19780 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 17296 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 22172 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 11776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 10212 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 9200 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 19596 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 9108 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 21988 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 18584 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 9384 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold41
timestamp 1679235063
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 21068 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold44
timestamp 1679235063
transform 1 0 10856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 9384 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 8280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 22264 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 24564 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 10120 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 24564 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 16376 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 15640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 5704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 4600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold61
timestamp 1679235063
transform 1 0 6900 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 14996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 6532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold65
timestamp 1679235063
transform 1 0 24380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 19504 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold68
timestamp 1679235063
transform 1 0 18032 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 6624 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1679235063
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 4416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform 1 0 20792 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold78
timestamp 1679235063
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform 1 0 6808 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold80
timestamp 1679235063
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold81
timestamp 1679235063
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold82
timestamp 1679235063
transform 1 0 16928 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 7636 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 23552 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform 1 0 6808 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1679235063
transform 1 0 11224 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold88
timestamp 1679235063
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold91
timestamp 1679235063
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold92
timestamp 1679235063
transform 1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold93
timestamp 1679235063
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 10948 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95
timestamp 1679235063
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform 1 0 11868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 14536 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 6808 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold99
timestamp 1679235063
transform 1 0 20424 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold100
timestamp 1679235063
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1679235063
transform 1 0 16836 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold102
timestamp 1679235063
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1679235063
transform 1 0 12236 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold105
timestamp 1679235063
transform 1 0 18216 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold106
timestamp 1679235063
transform 1 0 17940 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold107
timestamp 1679235063
transform 1 0 14628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold108
timestamp 1679235063
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold109
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1679235063
transform 1 0 9384 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold111
timestamp 1679235063
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold112
timestamp 1679235063
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold113
timestamp 1679235063
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold114
timestamp 1679235063
transform 1 0 17204 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold115
timestamp 1679235063
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold116
timestamp 1679235063
transform 1 0 7176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold117
timestamp 1679235063
transform 1 0 9292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold118
timestamp 1679235063
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold119
timestamp 1679235063
transform 1 0 5704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold120
timestamp 1679235063
transform 1 0 5612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold121
timestamp 1679235063
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold122
timestamp 1679235063
transform 1 0 6900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold123
timestamp 1679235063
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold124
timestamp 1679235063
transform 1 0 6716 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold125
timestamp 1679235063
transform 1 0 6532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold126
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold127
timestamp 1679235063
transform 1 0 2760 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold128
timestamp 1679235063
transform 1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold129
timestamp 1679235063
transform 1 0 24656 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold130
timestamp 1679235063
transform 1 0 24564 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold131
timestamp 1679235063
transform 1 0 22908 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold132
timestamp 1679235063
transform 1 0 22632 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold133
timestamp 1679235063
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold134
timestamp 1679235063
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold135
timestamp 1679235063
transform 1 0 23092 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold136
timestamp 1679235063
transform 1 0 24564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold137
timestamp 1679235063
transform 1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold138
timestamp 1679235063
transform 1 0 24196 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold139
timestamp 1679235063
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold140
timestamp 1679235063
transform 1 0 7176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold141
timestamp 1679235063
transform 1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold142
timestamp 1679235063
transform 1 0 8280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold143
timestamp 1679235063
transform 1 0 18032 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold144
timestamp 1679235063
transform 1 0 19412 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold145
timestamp 1679235063
transform 1 0 10856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold146
timestamp 1679235063
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold147
timestamp 1679235063
transform 1 0 17756 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold148
timestamp 1679235063
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold149
timestamp 1679235063
transform 1 0 19412 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold150
timestamp 1679235063
transform 1 0 23184 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold151
timestamp 1679235063
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold152
timestamp 1679235063
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold153
timestamp 1679235063
transform 1 0 15916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold154
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold155
timestamp 1679235063
transform 1 0 19596 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold156
timestamp 1679235063
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold157
timestamp 1679235063
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold158
timestamp 1679235063
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold159
timestamp 1679235063
transform 1 0 11684 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold160
timestamp 1679235063
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold161
timestamp 1679235063
transform 1 0 14720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold162
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold163
timestamp 1679235063
transform 1 0 11684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold164
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold165
timestamp 1679235063
transform 1 0 21988 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold166
timestamp 1679235063
transform 1 0 24380 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold167
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold168
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold169
timestamp 1679235063
transform 1 0 21528 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold170
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold171
timestamp 1679235063
transform 1 0 11684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold172
timestamp 1679235063
transform 1 0 12788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold173
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold174
timestamp 1679235063
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold175
timestamp 1679235063
transform 1 0 20240 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold176
timestamp 1679235063
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold177
timestamp 1679235063
transform 1 0 24564 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold178
timestamp 1679235063
transform 1 0 24564 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold179
timestamp 1679235063
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold180
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold181
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold182
timestamp 1679235063
transform 1 0 8280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold183
timestamp 1679235063
transform 1 0 18032 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold184
timestamp 1679235063
transform 1 0 18400 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold185
timestamp 1679235063
transform 1 0 17020 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold186
timestamp 1679235063
transform 1 0 23184 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold187
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold188
timestamp 1679235063
transform 1 0 11960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold189
timestamp 1679235063
transform 1 0 18492 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold190
timestamp 1679235063
transform 1 0 20700 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold191
timestamp 1679235063
transform 1 0 9936 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold192
timestamp 1679235063
transform 1 0 11316 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold193
timestamp 1679235063
transform 1 0 9016 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold194
timestamp 1679235063
transform 1 0 9752 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold195
timestamp 1679235063
transform 1 0 17940 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold196
timestamp 1679235063
transform 1 0 20700 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold197
timestamp 1679235063
transform 1 0 9752 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold198
timestamp 1679235063
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold199
timestamp 1679235063
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold200
timestamp 1679235063
transform 1 0 11684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold201
timestamp 1679235063
transform 1 0 19596 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold202
timestamp 1679235063
transform 1 0 22724 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold203
timestamp 1679235063
transform 1 0 24380 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold204
timestamp 1679235063
transform 1 0 6808 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold205
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold206
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold207
timestamp 1679235063
transform 1 0 15088 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold208
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold209
timestamp 1679235063
transform 1 0 17020 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold210
timestamp 1679235063
transform 1 0 18952 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold211
timestamp 1679235063
transform 1 0 11960 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold212
timestamp 1679235063
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold213
timestamp 1679235063
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold214
timestamp 1679235063
transform 1 0 24288 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold215
timestamp 1679235063
transform 1 0 9108 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold216
timestamp 1679235063
transform 1 0 9108 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold217
timestamp 1679235063
transform 1 0 20884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold218
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold219
timestamp 1679235063
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold220
timestamp 1679235063
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold221
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold222
timestamp 1679235063
transform 1 0 19044 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold223
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold224
timestamp 1679235063
transform 1 0 15732 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold225
timestamp 1679235063
transform 1 0 17940 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold226
timestamp 1679235063
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold227
timestamp 1679235063
transform 1 0 24656 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold228
timestamp 1679235063
transform 1 0 24564 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold229
timestamp 1679235063
transform 1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold230
timestamp 1679235063
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold231
timestamp 1679235063
transform 1 0 6900 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold232
timestamp 1679235063
transform 1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold233
timestamp 1679235063
transform 1 0 6808 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold234
timestamp 1679235063
transform 1 0 6808 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold235
timestamp 1679235063
transform 1 0 18216 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold236
timestamp 1679235063
transform 1 0 18400 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold237
timestamp 1679235063
transform 1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold238
timestamp 1679235063
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold239
timestamp 1679235063
transform 1 0 11684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold240
timestamp 1679235063
transform 1 0 11960 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold241
timestamp 1679235063
transform 1 0 24564 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold242
timestamp 1679235063
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold243
timestamp 1679235063
transform 1 0 4232 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1679235063
transform 1 0 4232 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold245
timestamp 1679235063
transform 1 0 5704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold246
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold247
timestamp 1679235063
transform 1 0 9384 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold248
timestamp 1679235063
transform 1 0 9476 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold249
timestamp 1679235063
transform 1 0 5152 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold250
timestamp 1679235063
transform 1 0 24656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold251
timestamp 1679235063
transform 1 0 19504 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold252
timestamp 1679235063
transform 1 0 20608 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold253
timestamp 1679235063
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1679235063
transform 1 0 4600 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold255
timestamp 1679235063
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold256
timestamp 1679235063
transform 1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold257
timestamp 1679235063
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold258
timestamp 1679235063
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold259
timestamp 1679235063
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1679235063
transform 1 0 3128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold261
timestamp 1679235063
transform 1 0 6808 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold262
timestamp 1679235063
transform 1 0 7544 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold263
timestamp 1679235063
transform 1 0 17112 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold264
timestamp 1679235063
transform 1 0 19596 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold265
timestamp 1679235063
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold266
timestamp 1679235063
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold267
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold268
timestamp 1679235063
transform 1 0 6808 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold269
timestamp 1679235063
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold270
timestamp 1679235063
transform 1 0 7912 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold271
timestamp 1679235063
transform 1 0 7728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold272
timestamp 1679235063
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold273
timestamp 1679235063
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold274
timestamp 1679235063
transform 1 0 7176 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold275
timestamp 1679235063
transform 1 0 24656 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold276
timestamp 1679235063
transform 1 0 24564 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold277
timestamp 1679235063
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold278
timestamp 1679235063
transform 1 0 6808 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold279
timestamp 1679235063
transform 1 0 16836 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold280
timestamp 1679235063
transform 1 0 15180 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold281
timestamp 1679235063
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold282
timestamp 1679235063
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold283
timestamp 1679235063
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold284
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold285
timestamp 1679235063
transform 1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold286
timestamp 1679235063
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold287
timestamp 1679235063
transform 1 0 4232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold288
timestamp 1679235063
transform 1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold289
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold290
timestamp 1679235063
transform 1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold291
timestamp 1679235063
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold292
timestamp 1679235063
transform 1 0 14444 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold293
timestamp 1679235063
transform 1 0 21528 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold294
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold295
timestamp 1679235063
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold296
timestamp 1679235063
transform 1 0 5704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold297
timestamp 1679235063
transform 1 0 24012 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold298
timestamp 1679235063
transform 1 0 22264 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold299
timestamp 1679235063
transform 1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold300
timestamp 1679235063
transform 1 0 6808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold301
timestamp 1679235063
transform 1 0 12788 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold302
timestamp 1679235063
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold303
timestamp 1679235063
transform 1 0 24656 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold304
timestamp 1679235063
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold305
timestamp 1679235063
transform 1 0 4232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold306
timestamp 1679235063
transform 1 0 11684 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold307
timestamp 1679235063
transform 1 0 12880 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold308
timestamp 1679235063
transform 1 0 8188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold309
timestamp 1679235063
transform 1 0 14628 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold310
timestamp 1679235063
transform 1 0 11684 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold311
timestamp 1679235063
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold312
timestamp 1679235063
transform 1 0 12880 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold313
timestamp 1679235063
transform 1 0 14536 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold314
timestamp 1679235063
transform 1 0 23184 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold315
timestamp 1679235063
transform 1 0 16836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold316
timestamp 1679235063
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold317
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold318
timestamp 1679235063
transform 1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold319
timestamp 1679235063
transform 1 0 7176 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold320
timestamp 1679235063
transform 1 0 9844 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold321
timestamp 1679235063
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold322
timestamp 1679235063
transform 1 0 10580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold323
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold324
timestamp 1679235063
transform 1 0 17112 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold325
timestamp 1679235063
transform 1 0 13340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold326
timestamp 1679235063
transform 1 0 17020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold327
timestamp 1679235063
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold328
timestamp 1679235063
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold329
timestamp 1679235063
transform 1 0 19412 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold330
timestamp 1679235063
transform 1 0 6716 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold331
timestamp 1679235063
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold332
timestamp 1679235063
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold333
timestamp 1679235063
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold334
timestamp 1679235063
transform 1 0 6808 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold335
timestamp 1679235063
transform 1 0 6808 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold336
timestamp 1679235063
transform 1 0 6808 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold337
timestamp 1679235063
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold338
timestamp 1679235063
transform 1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold339
timestamp 1679235063
transform 1 0 2668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold340
timestamp 1679235063
transform 1 0 3956 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold341
timestamp 1679235063
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold342
timestamp 1679235063
transform 1 0 3956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold343
timestamp 1679235063
transform 1 0 23460 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold344
timestamp 1679235063
transform 1 0 22264 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold345
timestamp 1679235063
transform 1 0 23368 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold346
timestamp 1679235063
transform 1 0 24564 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold347
timestamp 1679235063
transform 1 0 23092 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 23092 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 24012 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 23828 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1679235063
transform 1 0 22724 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1679235063
transform 1 0 25024 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1679235063
transform 1 0 25024 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 24380 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 24472 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1679235063
transform 1 0 25024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 12420 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1679235063
transform 1 0 25024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1679235063
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1679235063
transform 1 0 25024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 25116 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1679235063
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1679235063
transform 1 0 25024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1679235063
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 14352 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 23828 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 22080 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 21620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 18676 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 17848 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1679235063
transform 1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1679235063
transform 1 0 2576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1679235063
transform 1 0 7728 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1679235063
transform 1 0 2576 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1679235063
transform 1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1679235063
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1679235063
transform 1 0 1840 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1679235063
transform 1 0 3128 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1679235063
transform 1 0 3588 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1679235063
transform 1 0 2576 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1679235063
transform 1 0 2576 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1679235063
transform 1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1679235063
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform 1 0 4876 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1679235063
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 13524 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform 1 0 14904 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform 1 0 16836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 17664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1679235063
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input69
timestamp 1679235063
transform 1 0 24840 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1679235063
transform 1 0 24840 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1679235063
transform 1 0 24840 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24104 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1679235063
transform 1 0 21160 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1679235063
transform 1 0 22724 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1679235063
transform 1 0 22356 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform 1 0 23736 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 1564 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 17480 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 22080 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 20792 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 20056 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 12144 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 17296 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 17388 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 21988 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 19228 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 21620 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 23828 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 21252 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 20792 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 20056 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 17480 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 3956 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 5244 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 6624 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1679235063
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1679235063
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1679235063
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1679235063
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1679235063
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1679235063
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1679235063
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1679235063
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1679235063
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1679235063
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1679235063
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1679235063
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1679235063
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1679235063
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1679235063
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1679235063
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1679235063
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1679235063
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1679235063
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1679235063
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1679235063
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1679235063
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1679235063
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1679235063
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1679235063
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1679235063
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1679235063
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1679235063
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1679235063
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1679235063
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1679235063
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1679235063
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1679235063
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1679235063
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1679235063
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1679235063
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1679235063
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1679235063
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1679235063
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1679235063
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1679235063
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1679235063
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1679235063
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1679235063
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1679235063
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1679235063
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1679235063
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1679235063
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1679235063
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1679235063
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1679235063
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1679235063
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1679235063
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1679235063
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1679235063
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1679235063
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1679235063
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1679235063
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1679235063
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1679235063
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1679235063
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1679235063
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18400 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21436 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19044 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23092 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18032 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17572 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17020 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17664 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21068 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22724 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23368 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23368 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20608 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20516 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9844 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11040 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11224 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9384 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12604 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13064 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11776 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13984 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12788 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11316 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9384 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8556 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8556 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7268 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9660 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11592 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13984 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12880 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8832 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8740 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10580 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13984 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14076 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16284 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13432 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13064 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13984 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16008 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17848 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19872 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20608 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20424 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20332 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22172 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23000 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20424 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18216 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18216 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19596 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__201
timestamp 1679235063
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20148 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24196 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21436 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__165
timestamp 1679235063
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22356 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__166
timestamp 1679235063
transform 1 0 7268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__202
timestamp 1679235063
transform 1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__203
timestamp 1679235063
transform 1 0 9200 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4048 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__204
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19872 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22172 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18492 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__205
timestamp 1679235063
transform 1 0 20148 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 21620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20240 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 16928 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__157
timestamp 1679235063
transform 1 0 16468 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19596 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24196 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__159
timestamp 1679235063
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__160
timestamp 1679235063
transform 1 0 24932 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4324 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 19596 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__162
timestamp 1679235063
transform 1 0 19136 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19044 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23184 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22448 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__164
timestamp 1679235063
transform 1 0 2760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4416 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15364 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16560 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9568 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__167
timestamp 1679235063
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12052 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15456 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15456 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10212 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__173
timestamp 1679235063
transform 1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15916 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14812 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__184
timestamp 1679235063
transform 1 0 10948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14444 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16652 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17204 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10764 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__195
timestamp 1679235063
transform 1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11776 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14720 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16008 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12788 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__196
timestamp 1679235063
transform 1 0 6624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17940 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13984 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14444 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7084 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__168
timestamp 1679235063
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9568 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13524 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7820 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__169
timestamp 1679235063
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__170
timestamp 1679235063
transform 1 0 13432 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12880 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15916 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__171
timestamp 1679235063
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13800 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__172
timestamp 1679235063
transform 1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__174
timestamp 1679235063
transform 1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10488 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12328 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__175
timestamp 1679235063
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__176
timestamp 1679235063
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__177
timestamp 1679235063
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__178
timestamp 1679235063
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16008 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3772 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__179
timestamp 1679235063
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15272 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17572 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__180
timestamp 1679235063
transform 1 0 9476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18032 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16744 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12236 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__181
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16008 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 13248 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__182
timestamp 1679235063
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__183
timestamp 1679235063
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__185
timestamp 1679235063
transform 1 0 5060 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__186
timestamp 1679235063
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__187
timestamp 1679235063
transform 1 0 4416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18032 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19688 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2576 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__188
timestamp 1679235063
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__189
timestamp 1679235063
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__190
timestamp 1679235063
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__191
timestamp 1679235063
transform 1 0 5060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__192
timestamp 1679235063
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17756 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__193
timestamp 1679235063
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__194
timestamp 1679235063
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1679235063
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1679235063
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1679235063
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1679235063
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1679235063
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1679235063
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1679235063
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1679235063
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1679235063
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1679235063
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1679235063
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1679235063
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1679235063
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1679235063
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1679235063
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1679235063
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1679235063
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1679235063
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1679235063
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1679235063
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1679235063
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1679235063
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1679235063
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1679235063
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1679235063
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1679235063
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1679235063
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1679235063
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1679235063
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1679235063
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1679235063
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1679235063
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1679235063
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1679235063
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1679235063
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1679235063
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1679235063
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1679235063
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1679235063
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1679235063
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1679235063
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1679235063
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1679235063
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1679235063
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1679235063
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1679235063
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1679235063
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1679235063
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1679235063
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1679235063
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1679235063
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1679235063
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1679235063
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1679235063
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1679235063
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1679235063
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1679235063
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1679235063
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1679235063
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1679235063
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1679235063
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1679235063
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1679235063
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1679235063
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1679235063
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1679235063
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1679235063
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1679235063
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal2 10258 29410 10258 29410 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9982 45934 9982 45934 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9200 45390 9200 45390 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 8786 47532 8786 47532 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8188 39066 8188 39066 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 7958 16762 7958 16762 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 14582 8364 14582 8364 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 10902 13770 10902 13770 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 8464 13838 8464 13838 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 8924 15606 8924 15606 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 13386 13804 13386 13804 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 9246 10710 9246 10710 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal2 9798 13498 9798 13498 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal2 9660 23630 9660 23630 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal2 7774 16150 7774 16150 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal2 13616 19516 13616 19516 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 9752 18394 9752 18394 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 9706 20366 9706 20366 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 15594 18258 15594 18258 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 10810 24242 10810 24242 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 13984 8602 13984 8602 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9016 16422 9016 16422 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8648 32878 8648 32878 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12190 10608 12190 10608 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14582 9656 14582 9656 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 11960 12444 11960 12444 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10718 13226 10718 13226 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10626 15334 10626 15334 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11132 13940 11132 13940 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9200 13498 9200 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10258 14042 10258 14042 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9798 15572 9798 15572 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15502 7990 15502 7990 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9200 13770 9200 13770 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8832 17306 8832 17306 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15548 8330 15548 8330 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14214 9146 14214 9146 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15272 13158 15272 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12834 14008 12834 14008 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10810 11866 10810 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12604 10982 12604 10982 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9660 13770 9660 13770 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9568 14042 9568 14042 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10166 13498 10166 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14720 13294 14720 13294 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9936 23698 9936 23698 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9062 35666 9062 35666 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14582 10506 14582 10506 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13524 14314 13524 14314 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12788 14314 12788 14314 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12420 16218 12420 16218 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12972 13158 12972 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12650 15844 12650 15844 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10580 16218 10580 16218 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14674 21862 14674 21862 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9844 23834 9844 23834 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13984 16694 13984 16694 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10074 25299 10074 25299 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8832 38930 8832 38930 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14168 12410 14168 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 14909 12558 14909 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12650 12954 12650 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12926 17850 12926 17850 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12742 17697 12742 17697 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11730 15674 11730 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10488 18394 10488 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10442 24276 10442 24276 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10304 28390 10304 28390 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 11776 37842 11776 37842 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 10810 48994 10810 48994 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 15042 46002 15042 46002 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 9982 43146 9982 43146 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel via1 9522 45533 9522 45533 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 14674 47022 14674 47022 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 10534 45050 10534 45050 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 8878 50388 8878 50388 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 14490 47464 14490 47464 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5198 53040 5198 53040 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 11914 46614 11914 46614 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25070 53686 25070 53686 0 ccff_head
rlabel metal2 1518 1639 1518 1639 0 ccff_head_0
rlabel metal3 25676 748 25676 748 0 ccff_tail
rlabel metal1 1564 53618 1564 53618 0 ccff_tail_0
rlabel metal1 15364 26486 15364 26486 0 chanx_right_in[0]
rlabel metal1 24380 38930 24380 38930 0 chanx_right_in[10]
rlabel metal1 23138 38182 23138 38182 0 chanx_right_in[11]
rlabel metal1 23874 37706 23874 37706 0 chanx_right_in[12]
rlabel metal1 24748 39338 24748 39338 0 chanx_right_in[13]
rlabel metal1 24978 40086 24978 40086 0 chanx_right_in[14]
rlabel metal2 24702 39321 24702 39321 0 chanx_right_in[15]
rlabel metal2 25346 40103 25346 40103 0 chanx_right_in[16]
rlabel metal1 24748 40018 24748 40018 0 chanx_right_in[17]
rlabel metal1 24794 41106 24794 41106 0 chanx_right_in[18]
rlabel via2 25162 41531 25162 41531 0 chanx_right_in[19]
rlabel metal1 12305 27370 12305 27370 0 chanx_right_in[1]
rlabel metal2 25162 42483 25162 42483 0 chanx_right_in[20]
rlabel metal2 25530 43401 25530 43401 0 chanx_right_in[21]
rlabel metal2 24794 44183 24794 44183 0 chanx_right_in[22]
rlabel via2 25346 44829 25346 44829 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47447 25346 47447 0 chanx_right_in[26]
rlabel via2 25162 48093 25162 48093 0 chanx_right_in[27]
rlabel metal2 25162 49011 25162 49011 0 chanx_right_in[28]
rlabel metal2 25530 49929 25530 49929 0 chanx_right_in[29]
rlabel metal1 16744 29546 16744 29546 0 chanx_right_in[2]
rlabel metal1 24104 34918 24104 34918 0 chanx_right_in[3]
rlabel metal1 13800 29614 13800 29614 0 chanx_right_in[4]
rlabel metal1 23598 34918 23598 34918 0 chanx_right_in[5]
rlabel metal1 21942 32878 21942 32878 0 chanx_right_in[6]
rlabel metal2 22126 32419 22126 32419 0 chanx_right_in[7]
rlabel metal1 19458 35020 19458 35020 0 chanx_right_in[8]
rlabel metal2 22126 33915 22126 33915 0 chanx_right_in[9]
rlabel metal1 20700 2618 20700 2618 0 chanx_right_out[0]
rlabel metal2 25162 9129 25162 9129 0 chanx_right_out[10]
rlabel metal2 24794 10013 24794 10013 0 chanx_right_out[11]
rlabel metal1 24380 11050 24380 11050 0 chanx_right_out[12]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[13]
rlabel metal3 25584 12988 25584 12988 0 chanx_right_out[14]
rlabel metal1 23920 13362 23920 13362 0 chanx_right_out[15]
rlabel metal2 23322 15317 23322 15317 0 chanx_right_out[16]
rlabel metal3 25722 15436 25722 15436 0 chanx_right_out[17]
rlabel metal3 25722 16252 25722 16252 0 chanx_right_out[18]
rlabel metal2 25162 16609 25162 16609 0 chanx_right_out[19]
rlabel metal2 22218 2091 22218 2091 0 chanx_right_out[1]
rlabel metal1 24380 17714 24380 17714 0 chanx_right_out[20]
rlabel metal2 24794 17901 24794 17901 0 chanx_right_out[21]
rlabel metal2 23414 19635 23414 19635 0 chanx_right_out[22]
rlabel metal1 24426 19890 24426 19890 0 chanx_right_out[23]
rlabel via2 22494 21437 22494 21437 0 chanx_right_out[24]
rlabel metal1 24472 20978 24472 20978 0 chanx_right_out[25]
rlabel metal1 24012 22542 24012 22542 0 chanx_right_out[26]
rlabel metal1 24196 23154 24196 23154 0 chanx_right_out[27]
rlabel metal2 24794 23477 24794 23477 0 chanx_right_out[28]
rlabel metal3 25676 25228 25676 25228 0 chanx_right_out[29]
rlabel metal2 22310 6341 22310 6341 0 chanx_right_out[2]
rlabel metal1 13386 3128 13386 3128 0 chanx_right_out[3]
rlabel metal2 23322 8313 23322 8313 0 chanx_right_out[4]
rlabel metal2 24794 5389 24794 5389 0 chanx_right_out[5]
rlabel metal3 25722 6460 25722 6460 0 chanx_right_out[6]
rlabel metal2 24794 6749 24794 6749 0 chanx_right_out[7]
rlabel metal1 24380 7922 24380 7922 0 chanx_right_out[8]
rlabel metal1 24104 8398 24104 8398 0 chanx_right_out[9]
rlabel metal2 1886 823 1886 823 0 chany_bottom_in_0[0]
rlabel metal1 1334 12614 1334 12614 0 chany_bottom_in_0[10]
rlabel metal2 5934 823 5934 823 0 chany_bottom_in_0[11]
rlabel metal1 4462 9690 4462 9690 0 chany_bottom_in_0[12]
rlabel metal1 4002 10540 4002 10540 0 chany_bottom_in_0[13]
rlabel metal2 2714 11390 2714 11390 0 chany_bottom_in_0[14]
rlabel metal2 1978 11628 1978 11628 0 chany_bottom_in_0[15]
rlabel metal2 874 9146 874 9146 0 chany_bottom_in_0[16]
rlabel metal1 2346 6766 2346 6766 0 chany_bottom_in_0[17]
rlabel metal2 2070 14297 2070 14297 0 chany_bottom_in_0[18]
rlabel metal1 1610 10030 1610 10030 0 chany_bottom_in_0[19]
rlabel metal1 1840 9554 1840 9554 0 chany_bottom_in_0[1]
rlabel via2 3818 12597 3818 12597 0 chany_bottom_in_0[20]
rlabel metal1 1380 15402 1380 15402 0 chany_bottom_in_0[21]
rlabel metal1 1886 6154 1886 6154 0 chany_bottom_in_0[22]
rlabel metal1 1702 14858 1702 14858 0 chany_bottom_in_0[23]
rlabel metal1 1702 15470 1702 15470 0 chany_bottom_in_0[24]
rlabel metal1 3634 15402 3634 15402 0 chany_bottom_in_0[25]
rlabel metal2 11730 3196 11730 3196 0 chany_bottom_in_0[26]
rlabel metal2 3404 2516 3404 2516 0 chany_bottom_in_0[27]
rlabel metal2 12190 1367 12190 1367 0 chany_bottom_in_0[28]
rlabel metal2 12466 527 12466 527 0 chany_bottom_in_0[29]
rlabel metal1 2622 3604 2622 3604 0 chany_bottom_in_0[2]
rlabel metal2 2944 2516 2944 2516 0 chany_bottom_in_0[3]
rlabel metal1 3174 2482 3174 2482 0 chany_bottom_in_0[4]
rlabel metal2 3726 1095 3726 1095 0 chany_bottom_in_0[5]
rlabel metal2 4094 1095 4094 1095 0 chany_bottom_in_0[6]
rlabel metal2 2070 11339 2070 11339 0 chany_bottom_in_0[7]
rlabel metal2 6532 14994 6532 14994 0 chany_bottom_in_0[8]
rlabel metal1 5520 2414 5520 2414 0 chany_bottom_in_0[9]
rlabel metal2 12926 1231 12926 1231 0 chany_bottom_out_0[0]
rlabel metal2 16606 959 16606 959 0 chany_bottom_out_0[10]
rlabel metal1 17710 3638 17710 3638 0 chany_bottom_out_0[11]
rlabel metal1 17848 3706 17848 3706 0 chany_bottom_out_0[12]
rlabel metal2 17710 1690 17710 1690 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal2 18446 1707 18446 1707 0 chany_bottom_out_0[15]
rlabel metal1 19780 3162 19780 3162 0 chany_bottom_out_0[16]
rlabel metal2 19182 1761 19182 1761 0 chany_bottom_out_0[17]
rlabel metal1 20516 2958 20516 2958 0 chany_bottom_out_0[18]
rlabel metal2 19918 1792 19918 1792 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal1 20930 4114 20930 4114 0 chany_bottom_out_0[20]
rlabel metal2 20654 1761 20654 1761 0 chany_bottom_out_0[21]
rlabel metal2 21022 1571 21022 1571 0 chany_bottom_out_0[22]
rlabel metal2 21390 2370 21390 2370 0 chany_bottom_out_0[23]
rlabel metal2 21758 3492 21758 3492 0 chany_bottom_out_0[24]
rlabel metal2 21942 5015 21942 5015 0 chany_bottom_out_0[25]
rlabel metal1 22264 7786 22264 7786 0 chany_bottom_out_0[26]
rlabel metal2 22862 1761 22862 1761 0 chany_bottom_out_0[27]
rlabel metal2 23230 1690 23230 1690 0 chany_bottom_out_0[28]
rlabel metal1 21850 5746 21850 5746 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14398 3570 14398 3570 0 chany_bottom_out_0[3]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal2 15134 1622 15134 1622 0 chany_bottom_out_0[6]
rlabel metal1 16054 3570 16054 3570 0 chany_bottom_out_0[7]
rlabel metal1 16606 2958 16606 2958 0 chany_bottom_out_0[8]
rlabel metal1 17710 2890 17710 2890 0 chany_bottom_out_0[9]
rlabel metal2 19734 16660 19734 16660 0 clknet_0_prog_clk
rlabel metal2 9430 13430 9430 13430 0 clknet_4_0_0_prog_clk
rlabel metal1 11638 42534 11638 42534 0 clknet_4_10_0_prog_clk
rlabel metal2 12650 29648 12650 29648 0 clknet_4_11_0_prog_clk
rlabel metal1 17618 26962 17618 26962 0 clknet_4_12_0_prog_clk
rlabel metal1 21988 24174 21988 24174 0 clknet_4_13_0_prog_clk
rlabel metal2 19458 32436 19458 32436 0 clknet_4_14_0_prog_clk
rlabel metal1 20010 43758 20010 43758 0 clknet_4_15_0_prog_clk
rlabel metal1 13064 5134 13064 5134 0 clknet_4_1_0_prog_clk
rlabel metal2 7268 22100 7268 22100 0 clknet_4_2_0_prog_clk
rlabel metal1 13938 19346 13938 19346 0 clknet_4_3_0_prog_clk
rlabel metal1 17710 12614 17710 12614 0 clknet_4_4_0_prog_clk
rlabel metal2 22034 8160 22034 8160 0 clknet_4_5_0_prog_clk
rlabel metal1 16928 20434 16928 20434 0 clknet_4_6_0_prog_clk
rlabel metal1 19734 19414 19734 19414 0 clknet_4_7_0_prog_clk
rlabel metal1 11822 27948 11822 27948 0 clknet_4_8_0_prog_clk
rlabel metal1 11178 25330 11178 25330 0 clknet_4_9_0_prog_clk
rlabel metal1 2484 54094 2484 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 4002 56236 4002 56236 0 gfpga_pad_io_soc_dir[1]
rlabel metal1 5474 53618 5474 53618 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6762 56236 6762 56236 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 13616 54162 13616 54162 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14996 54162 14996 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16836 54162 16836 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 17756 54162 17756 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal2 9338 51894 9338 51894 0 gfpga_pad_io_soc_out[1]
rlabel metal2 10902 56236 10902 56236 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12098 51112 12098 51112 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54094 19228 54094 0 isol_n
rlabel metal1 23230 52666 23230 52666 0 net1
rlabel metal2 24932 38420 24932 38420 0 net10
rlabel metal1 22632 25262 22632 25262 0 net100
rlabel metal2 17066 1088 17066 1088 0 net101
rlabel metal2 12190 4692 12190 4692 0 net102
rlabel metal2 12834 8211 12834 8211 0 net103
rlabel via3 12029 18020 12029 18020 0 net104
rlabel via2 20102 6715 20102 6715 0 net105
rlabel metal4 15824 15980 15824 15980 0 net106
rlabel metal1 20930 7820 20930 7820 0 net107
rlabel metal3 18469 1972 18469 1972 0 net108
rlabel metal1 21252 12614 21252 12614 0 net109
rlabel metal1 24748 32946 24748 32946 0 net11
rlabel metal3 16583 15300 16583 15300 0 net110
rlabel metal2 14766 4981 14766 4981 0 net111
rlabel metal1 16882 5202 16882 5202 0 net112
rlabel metal1 21942 2414 21942 2414 0 net113
rlabel via3 14237 20740 14237 20740 0 net114
rlabel metal1 14812 4726 14812 4726 0 net115
rlabel metal3 15295 1836 15295 1836 0 net116
rlabel metal1 20424 5338 20424 5338 0 net117
rlabel metal1 16376 17578 16376 17578 0 net118
rlabel metal1 18630 18870 18630 18870 0 net119
rlabel metal1 24196 40902 24196 40902 0 net12
rlabel metal2 12558 2057 12558 2057 0 net120
rlabel metal2 2714 6018 2714 6018 0 net121
rlabel metal2 20746 6936 20746 6936 0 net122
rlabel via3 9821 16660 9821 16660 0 net123
rlabel metal2 15134 3383 15134 3383 0 net124
rlabel metal2 5106 5831 5106 5831 0 net125
rlabel metal1 2760 2618 2760 2618 0 net126
rlabel metal3 12788 6936 12788 6936 0 net127
rlabel metal2 16606 9469 16606 9469 0 net128
rlabel metal3 18630 8364 18630 8364 0 net129
rlabel metal2 24886 41497 24886 41497 0 net13
rlabel metal2 2162 3638 2162 3638 0 net130
rlabel metal1 17618 2550 17618 2550 0 net131
rlabel metal2 14490 3621 14490 3621 0 net132
rlabel metal1 17641 2278 17641 2278 0 net133
rlabel metal1 15824 3026 15824 3026 0 net134
rlabel metal1 17112 2414 17112 2414 0 net135
rlabel metal2 16238 5338 16238 5338 0 net136
rlabel metal1 15962 13430 15962 13430 0 net137
rlabel metal2 18906 5168 18906 5168 0 net138
rlabel metal1 4462 53210 4462 53210 0 net139
rlabel metal2 13754 27013 13754 27013 0 net14
rlabel metal2 6578 53686 6578 53686 0 net140
rlabel metal2 7682 53108 7682 53108 0 net141
rlabel metal2 6762 53142 6762 53142 0 net142
rlabel metal2 7774 14416 7774 14416 0 net143
rlabel metal1 1978 6834 1978 6834 0 net144
rlabel metal1 24288 2618 24288 2618 0 net145
rlabel via1 13393 16150 13393 16150 0 net146
rlabel metal1 14451 21590 14451 21590 0 net147
rlabel metal2 20102 14756 20102 14756 0 net148
rlabel metal2 18998 21284 18998 21284 0 net149
rlabel metal2 25254 42585 25254 42585 0 net15
rlabel metal1 21397 26350 21397 26350 0 net150
rlabel metal1 22349 33898 22349 33898 0 net151
rlabel via1 11822 28475 11822 28475 0 net152
rlabel metal1 21199 43690 21199 43690 0 net153
rlabel metal2 18446 26146 18446 26146 0 net154
rlabel metal2 16974 28322 16974 28322 0 net155
rlabel metal1 18860 16626 18860 16626 0 net156
rlabel metal1 18446 29274 18446 29274 0 net157
rlabel metal2 21942 27710 21942 27710 0 net158
rlabel metal1 23184 32538 23184 32538 0 net159
rlabel metal2 23506 41565 23506 41565 0 net16
rlabel metal1 23690 29206 23690 29206 0 net160
rlabel metal1 20286 30192 20286 30192 0 net161
rlabel metal2 19826 29886 19826 29886 0 net162
rlabel metal1 19182 18156 19182 18156 0 net163
rlabel metal1 22862 17136 22862 17136 0 net164
rlabel metal1 10994 24684 10994 24684 0 net165
rlabel metal1 8234 23222 8234 23222 0 net166
rlabel metal1 3266 17782 3266 17782 0 net167
rlabel metal1 5382 12886 5382 12886 0 net168
rlabel metal1 5750 12138 5750 12138 0 net169
rlabel metal1 19872 44234 19872 44234 0 net17
rlabel metal1 13386 18394 13386 18394 0 net170
rlabel metal1 15180 17238 15180 17238 0 net171
rlabel metal2 14674 16218 14674 16218 0 net172
rlabel metal1 10718 20570 10718 20570 0 net173
rlabel metal1 11408 10030 11408 10030 0 net174
rlabel metal2 12558 7208 12558 7208 0 net175
rlabel metal1 13202 5100 13202 5100 0 net176
rlabel metal1 11086 11866 11086 11866 0 net177
rlabel metal1 14950 14994 14950 14994 0 net178
rlabel metal1 15272 16218 15272 16218 0 net179
rlabel metal1 23782 44710 23782 44710 0 net18
rlabel metal2 9522 14926 9522 14926 0 net180
rlabel metal1 12098 2482 12098 2482 0 net181
rlabel metal3 11086 1428 11086 1428 0 net182
rlabel metal1 1748 14042 1748 14042 0 net183
rlabel metal1 11592 21522 11592 21522 0 net184
rlabel metal2 5382 2193 5382 2193 0 net185
rlabel metal2 21114 10115 21114 10115 0 net186
rlabel metal1 5290 11798 5290 11798 0 net187
rlabel via2 19366 13515 19366 13515 0 net188
rlabel metal1 19228 11186 19228 11186 0 net189
rlabel metal1 23828 45798 23828 45798 0 net19
rlabel via2 3266 9979 3266 9979 0 net190
rlabel metal2 20746 5151 20746 5151 0 net191
rlabel metal2 1702 6137 1702 6137 0 net192
rlabel metal3 1541 9724 1541 9724 0 net193
rlabel metal1 10672 7786 10672 7786 0 net194
rlabel metal1 5842 17748 5842 17748 0 net195
rlabel metal1 9016 17578 9016 17578 0 net196
rlabel metal1 5980 13838 5980 13838 0 net197
rlabel metal1 13570 9486 13570 9486 0 net198
rlabel metal1 14444 21998 14444 21998 0 net199
rlabel metal2 3910 9843 3910 9843 0 net2
rlabel metal1 23920 46342 23920 46342 0 net20
rlabel metal1 15962 23834 15962 23834 0 net200
rlabel metal2 24012 19244 24012 19244 0 net201
rlabel metal2 9154 22389 9154 22389 0 net202
rlabel metal1 9246 26418 9246 26418 0 net203
rlabel metal2 20286 23732 20286 23732 0 net204
rlabel metal1 20102 18394 20102 18394 0 net205
rlabel metal2 4002 6052 4002 6052 0 net206
rlabel metal2 4830 4284 4830 4284 0 net207
rlabel metal1 25208 53210 25208 53210 0 net208
rlabel metal2 22678 48042 22678 48042 0 net209
rlabel metal1 25484 47430 25484 47430 0 net21
rlabel metal1 20838 18224 20838 18224 0 net210
rlabel metal1 24932 26962 24932 26962 0 net211
rlabel metal2 24242 35326 24242 35326 0 net212
rlabel metal1 7084 3026 7084 3026 0 net213
rlabel metal1 10764 23834 10764 23834 0 net214
rlabel metal2 18630 26826 18630 26826 0 net215
rlabel metal1 12972 4590 12972 4590 0 net216
rlabel metal1 13248 5678 13248 5678 0 net217
rlabel metal1 22954 31450 22954 31450 0 net218
rlabel metal1 16376 15130 16376 15130 0 net219
rlabel metal3 22701 46988 22701 46988 0 net22
rlabel metal1 20516 34578 20516 34578 0 net220
rlabel metal1 18262 33626 18262 33626 0 net221
rlabel metal1 18262 5746 18262 5746 0 net222
rlabel metal2 24426 29852 24426 29852 0 net223
rlabel metal2 10534 27710 10534 27710 0 net224
rlabel metal2 13110 24004 13110 24004 0 net225
rlabel metal3 7797 1292 7797 1292 0 net226
rlabel metal1 25162 14246 25162 14246 0 net227
rlabel metal1 11408 20434 11408 20434 0 net228
rlabel metal1 20654 28186 20654 28186 0 net229
rlabel metal2 25254 48297 25254 48297 0 net23
rlabel metal2 25254 34612 25254 34612 0 net230
rlabel metal1 18262 12240 18262 12240 0 net231
rlabel metal1 8464 12818 8464 12818 0 net232
rlabel metal1 11500 30294 11500 30294 0 net233
rlabel metal1 24932 2618 24932 2618 0 net234
rlabel metal1 18216 31314 18216 31314 0 net235
rlabel metal1 23046 36006 23046 36006 0 net236
rlabel metal2 12466 8772 12466 8772 0 net237
rlabel metal2 10902 44676 10902 44676 0 net238
rlabel metal1 9844 31994 9844 31994 0 net239
rlabel metal3 22931 47668 22931 47668 0 net24
rlabel metal1 20516 35054 20516 35054 0 net240
rlabel metal1 9476 47226 9476 47226 0 net241
rlabel metal2 24610 24922 24610 24922 0 net242
rlabel metal2 19090 18700 19090 18700 0 net243
rlabel metal2 10074 3604 10074 3604 0 net244
rlabel metal1 11730 5644 11730 5644 0 net245
rlabel metal1 20286 23222 20286 23222 0 net246
rlabel metal2 20746 22780 20746 22780 0 net247
rlabel metal2 18998 9724 18998 9724 0 net248
rlabel metal2 10534 4284 10534 4284 0 net249
rlabel metal1 18584 20026 18584 20026 0 net25
rlabel metal1 10304 5202 10304 5202 0 net250
rlabel metal2 6854 26554 6854 26554 0 net251
rlabel metal1 24012 11322 24012 11322 0 net252
rlabel metal1 17204 22746 17204 22746 0 net253
rlabel metal1 23184 36550 23184 36550 0 net254
rlabel metal1 25070 31926 25070 31926 0 net255
rlabel metal1 11960 29138 11960 29138 0 net256
rlabel metal1 9200 6766 9200 6766 0 net257
rlabel metal2 25254 36788 25254 36788 0 net258
rlabel metal2 18446 14076 18446 14076 0 net259
rlabel metal1 24748 33830 24748 33830 0 net26
rlabel metal1 16928 20026 16928 20026 0 net260
rlabel metal1 15732 26554 15732 26554 0 net261
rlabel metal1 9200 5678 9200 5678 0 net262
rlabel metal1 5566 10098 5566 10098 0 net263
rlabel metal1 5704 14994 5704 14994 0 net264
rlabel metal3 14145 18020 14145 18020 0 net265
rlabel via2 7222 23613 7222 23613 0 net266
rlabel metal2 6026 18564 6026 18564 0 net267
rlabel metal1 18262 17102 18262 17102 0 net268
rlabel metal2 7222 8772 7222 8772 0 net269
rlabel metal2 21942 25364 21942 25364 0 net27
rlabel metal4 15180 19108 15180 19108 0 net270
rlabel metal1 20424 25874 20424 25874 0 net271
rlabel metal1 5704 7378 5704 7378 0 net272
rlabel metal3 17388 748 17388 748 0 net273
rlabel metal1 7728 21522 7728 21522 0 net274
rlabel metal2 7314 9826 7314 9826 0 net275
rlabel metal2 10534 9996 10534 9996 0 net276
rlabel metal2 15226 25534 15226 25534 0 net277
rlabel metal1 7912 3162 7912 3162 0 net278
rlabel metal1 5244 15674 5244 15674 0 net279
rlabel metal2 22724 34612 22724 34612 0 net28
rlabel metal2 5934 16864 5934 16864 0 net280
rlabel metal1 7774 5338 7774 5338 0 net281
rlabel metal1 20010 10642 20010 10642 0 net282
rlabel metal2 18906 14875 18906 14875 0 net283
rlabel metal2 6854 20876 6854 20876 0 net284
rlabel metal1 5474 12410 5474 12410 0 net285
rlabel metal1 22862 17272 22862 17272 0 net286
rlabel metal1 24472 19822 24472 19822 0 net287
rlabel metal2 8326 8772 8326 8772 0 net288
rlabel metal1 14720 11322 14720 11322 0 net289
rlabel metal2 21666 32368 21666 32368 0 net29
rlabel metal1 24426 36890 24426 36890 0 net290
rlabel metal1 6440 14314 6440 14314 0 net291
rlabel metal2 11914 41242 11914 41242 0 net292
rlabel metal1 7912 5882 7912 5882 0 net293
rlabel metal1 22310 37196 22310 37196 0 net294
rlabel metal2 12282 19176 12282 19176 0 net295
rlabel via2 6026 11645 6026 11645 0 net296
rlabel metal1 15686 31348 15686 31348 0 net297
rlabel metal1 9890 3910 9890 3910 0 net298
rlabel metal1 11592 26282 11592 26282 0 net299
rlabel metal3 18699 14756 18699 14756 0 net3
rlabel metal1 19090 33286 19090 33286 0 net30
rlabel metal2 13202 21726 13202 21726 0 net300
rlabel metal1 12512 27098 12512 27098 0 net301
rlabel metal1 14812 18394 14812 18394 0 net302
rlabel metal1 7590 11322 7590 11322 0 net303
rlabel metal1 21068 17850 21068 17850 0 net304
rlabel metal1 7721 13702 7721 13702 0 net305
rlabel metal1 14069 28934 14069 28934 0 net306
rlabel metal2 16146 15759 16146 15759 0 net307
rlabel metal1 10251 27642 10251 27642 0 net308
rlabel metal2 21298 14025 21298 14025 0 net309
rlabel metal2 22356 34068 22356 34068 0 net31
rlabel metal2 14582 35020 14582 35020 0 net310
rlabel metal2 18630 21250 18630 21250 0 net311
rlabel metal2 15318 21563 15318 21563 0 net312
rlabel metal1 8510 24718 8510 24718 0 net313
rlabel metal1 17020 13158 17020 13158 0 net314
rlabel metal1 9890 26758 9890 26758 0 net315
rlabel metal1 9752 29206 9752 29206 0 net316
rlabel metal1 11316 14994 11316 14994 0 net317
rlabel metal1 8786 26554 8786 26554 0 net318
rlabel metal2 17158 18462 17158 18462 0 net319
rlabel metal1 18906 34374 18906 34374 0 net32
rlabel metal1 6394 20570 6394 20570 0 net320
rlabel metal2 20930 1717 20930 1717 0 net321
rlabel metal1 9568 23018 9568 23018 0 net322
rlabel metal1 17480 10234 17480 10234 0 net323
rlabel metal1 6808 18666 6808 18666 0 net324
rlabel metal1 9880 20026 9880 20026 0 net325
rlabel metal1 10304 17714 10304 17714 0 net326
rlabel metal1 9006 14586 9006 14586 0 net327
rlabel metal1 6762 8058 6762 8058 0 net328
rlabel metal1 9476 10710 9476 10710 0 net329
rlabel metal1 11454 7922 11454 7922 0 net33
rlabel metal1 4830 2516 4830 2516 0 net330
rlabel metal1 3680 2550 3680 2550 0 net331
rlabel metal1 3726 4590 3726 4590 0 net332
rlabel metal1 5428 4250 5428 4250 0 net333
rlabel metal2 25346 53448 25346 53448 0 net334
rlabel metal2 25254 53958 25254 53958 0 net335
rlabel metal2 22586 50490 22586 50490 0 net336
rlabel metal1 22080 46954 22080 46954 0 net337
rlabel metal1 22034 18292 22034 18292 0 net338
rlabel metal2 22126 19958 22126 19958 0 net339
rlabel metal1 13340 14042 13340 14042 0 net34
rlabel metal1 24196 29614 24196 29614 0 net340
rlabel metal1 24472 27098 24472 27098 0 net341
rlabel metal1 20884 36142 20884 36142 0 net342
rlabel metal2 24886 34272 24886 34272 0 net343
rlabel metal1 6716 10626 6716 10626 0 net344
rlabel metal1 13754 986 13754 986 0 net345
rlabel metal1 10534 23664 10534 23664 0 net346
rlabel metal1 9190 25466 9190 25466 0 net347
rlabel metal2 18722 25908 18722 25908 0 net348
rlabel metal2 20102 27778 20102 27778 0 net349
rlabel metal1 12052 12206 12052 12206 0 net35
rlabel metal1 11776 3706 11776 3706 0 net350
rlabel metal1 14996 4522 14996 4522 0 net351
rlabel metal2 18446 33286 18446 33286 0 net352
rlabel metal1 18262 32334 18262 32334 0 net353
rlabel metal1 20562 30838 20562 30838 0 net354
rlabel metal1 20746 31892 20746 31892 0 net355
rlabel metal1 14398 6290 14398 6290 0 net356
rlabel metal2 13386 5406 13386 5406 0 net357
rlabel metal2 16606 14790 16606 14790 0 net358
rlabel metal1 16376 16150 16376 16150 0 net359
rlabel metal2 2622 8432 2622 8432 0 net36
rlabel metal2 19642 34748 19642 34748 0 net360
rlabel metal1 20562 34714 20562 34714 0 net361
rlabel metal1 16284 7446 16284 7446 0 net362
rlabel metal1 18170 5882 18170 5882 0 net363
rlabel metal1 11546 25806 11546 25806 0 net364
rlabel metal1 11270 27098 11270 27098 0 net365
rlabel metal1 13156 23698 13156 23698 0 net366
rlabel metal1 14720 24310 14720 24310 0 net367
rlabel metal1 11960 18394 11960 18394 0 net368
rlabel metal1 12144 20570 12144 20570 0 net369
rlabel metal2 2714 10285 2714 10285 0 net37
rlabel metal1 23000 30702 23000 30702 0 net370
rlabel metal2 23322 28322 23322 28322 0 net371
rlabel metal1 24886 14382 24886 14382 0 net372
rlabel metal1 25300 12410 25300 12410 0 net373
rlabel metal2 14582 18649 14582 18649 0 net374
rlabel metal1 24702 18190 24702 18190 0 net375
rlabel metal2 10534 31042 10534 31042 0 net376
rlabel metal2 12926 30430 12926 30430 0 net377
rlabel metal1 20056 10234 20056 10234 0 net378
rlabel metal1 18814 12410 18814 12410 0 net379
rlabel metal1 6210 12954 6210 12954 0 net38
rlabel metal2 20930 27574 20930 27574 0 net380
rlabel metal1 19458 29206 19458 29206 0 net381
rlabel metal1 25162 33966 25162 33966 0 net382
rlabel metal1 25116 34918 25116 34918 0 net383
rlabel metal2 24610 1972 24610 1972 0 net384
rlabel metal2 17342 6732 17342 6732 0 net385
rlabel metal1 11776 13906 11776 13906 0 net386
rlabel metal1 9338 12750 9338 12750 0 net387
rlabel metal1 18308 30294 18308 30294 0 net388
rlabel metal2 17434 30940 17434 30940 0 net389
rlabel metal1 9430 10540 9430 10540 0 net39
rlabel metal1 18814 33898 18814 33898 0 net390
rlabel metal2 20838 34476 20838 34476 0 net391
rlabel metal2 10718 8228 10718 8228 0 net392
rlabel metal2 12650 9316 12650 9316 0 net393
rlabel metal2 19182 35190 19182 35190 0 net394
rlabel metal1 20056 32946 20056 32946 0 net395
rlabel metal1 10442 43962 10442 43962 0 net396
rlabel metal1 11362 44778 11362 44778 0 net397
rlabel metal2 9706 31042 9706 31042 0 net398
rlabel metal1 10074 34170 10074 34170 0 net399
rlabel metal1 22586 38726 22586 38726 0 net4
rlabel metal1 14812 2346 14812 2346 0 net40
rlabel metal1 20884 23086 20884 23086 0 net400
rlabel metal2 21390 23732 21390 23732 0 net401
rlabel metal2 9430 3196 9430 3196 0 net402
rlabel metal2 18538 3485 18538 3485 0 net403
rlabel metal1 6854 6732 6854 6732 0 net404
rlabel metal1 11776 5882 11776 5882 0 net405
rlabel metal2 20286 11356 20286 11356 0 net406
rlabel metal1 22540 19278 22540 19278 0 net407
rlabel metal1 9246 27302 9246 27302 0 net408
rlabel metal1 10028 26418 10028 26418 0 net409
rlabel metal2 16238 13974 16238 13974 0 net41
rlabel metal2 20194 22780 20194 22780 0 net410
rlabel metal1 25622 16558 25622 16558 0 net411
rlabel metal1 16238 21658 16238 21658 0 net412
rlabel metal1 14904 22542 14904 22542 0 net413
rlabel metal1 17986 10030 17986 10030 0 net414
rlabel metal1 20286 15402 20286 15402 0 net415
rlabel metal1 10902 4556 10902 4556 0 net416
rlabel metal1 13386 4012 13386 4012 0 net417
rlabel metal1 23138 36346 23138 36346 0 net418
rlabel metal1 23138 33422 23138 33422 0 net419
rlabel metal2 1886 14093 1886 14093 0 net42
rlabel metal2 9798 46580 9798 46580 0 net420
rlabel metal1 6854 48008 6854 48008 0 net421
rlabel metal2 21574 25126 21574 25126 0 net422
rlabel metal1 25208 24378 25208 24378 0 net423
rlabel metal1 10580 3094 10580 3094 0 net424
rlabel metal1 13156 5338 13156 5338 0 net425
rlabel metal1 18860 19346 18860 19346 0 net426
rlabel metal1 19504 18394 19504 18394 0 net427
rlabel metal2 17526 19652 17526 19652 0 net428
rlabel metal1 15640 20366 15640 20366 0 net429
rlabel metal1 1610 10132 1610 10132 0 net43
rlabel metal1 16192 26350 16192 26350 0 net430
rlabel metal2 13754 27710 13754 27710 0 net431
rlabel metal2 24610 36346 24610 36346 0 net432
rlabel metal1 25346 37094 25346 37094 0 net433
rlabel metal2 6210 15878 6210 15878 0 net434
rlabel metal1 7176 14926 7176 14926 0 net435
rlabel metal1 5382 18224 5382 18224 0 net436
rlabel metal2 6026 19040 6026 19040 0 net437
rlabel metal2 7498 8262 7498 8262 0 net438
rlabel metal2 18722 8959 18722 8959 0 net439
rlabel metal1 1656 9418 1656 9418 0 net44
rlabel metal2 18262 14586 18262 14586 0 net440
rlabel metal2 19090 14790 19090 14790 0 net441
rlabel metal1 9844 4522 9844 4522 0 net442
rlabel metal1 13386 7344 13386 7344 0 net443
rlabel metal1 10166 29648 10166 29648 0 net444
rlabel metal2 11546 29410 11546 29410 0 net445
rlabel metal1 24932 31790 24932 31790 0 net446
rlabel metal1 23414 29750 23414 29750 0 net447
rlabel metal2 1518 8245 1518 8245 0 net448
rlabel metal3 18492 20536 18492 20536 0 net449
rlabel metal1 2622 12852 2622 12852 0 net45
rlabel metal2 6946 23868 6946 23868 0 net450
rlabel metal1 24702 13498 24702 13498 0 net451
rlabel metal1 7958 7888 7958 7888 0 net452
rlabel metal2 10166 7038 10166 7038 0 net453
rlabel metal2 4692 18292 4692 18292 0 net454
rlabel metal1 24886 18598 24886 18598 0 net455
rlabel metal1 19872 25466 19872 25466 0 net456
rlabel metal2 21298 26452 21298 26452 0 net457
rlabel metal2 5750 10234 5750 10234 0 net458
rlabel metal2 5474 8483 5474 8483 0 net459
rlabel metal1 17664 6086 17664 6086 0 net46
rlabel metal1 8878 11118 8878 11118 0 net460
rlabel metal1 10166 9146 10166 9146 0 net461
rlabel metal2 8326 3196 8326 3196 0 net462
rlabel metal1 13616 850 13616 850 0 net463
rlabel metal3 15180 4148 15180 4148 0 net464
rlabel via2 22034 14331 22034 14331 0 net465
rlabel metal1 5290 16524 5290 16524 0 net466
rlabel metal1 8280 16150 8280 16150 0 net467
rlabel metal1 19320 11118 19320 11118 0 net468
rlabel metal2 20286 10846 20286 10846 0 net469
rlabel metal2 2346 3961 2346 3961 0 net47
rlabel metal2 5382 8636 5382 8636 0 net470
rlabel metal2 6854 7463 6854 7463 0 net471
rlabel metal1 6854 21556 6854 21556 0 net472
rlabel metal1 8004 20366 8004 20366 0 net473
rlabel metal1 6854 24140 6854 24140 0 net474
rlabel metal1 8740 21658 8740 21658 0 net475
rlabel metal2 7682 8908 7682 8908 0 net476
rlabel metal1 8832 8534 8832 8534 0 net477
rlabel metal1 7774 5678 7774 5678 0 net478
rlabel metal1 8786 6358 8786 6358 0 net479
rlabel metal1 14950 8330 14950 8330 0 net48
rlabel metal1 23598 36788 23598 36788 0 net480
rlabel metal1 25116 38182 25116 38182 0 net481
rlabel metal1 6348 9554 6348 9554 0 net482
rlabel metal2 16422 9911 16422 9911 0 net483
rlabel metal2 16790 26554 16790 26554 0 net484
rlabel metal1 15686 24786 15686 24786 0 net485
rlabel metal1 4692 15130 4692 15130 0 net486
rlabel metal1 6578 16626 6578 16626 0 net487
rlabel metal1 20516 20570 20516 20570 0 net488
rlabel metal1 24058 20026 24058 20026 0 net489
rlabel metal2 19274 13124 19274 13124 0 net49
rlabel metal1 7176 5202 7176 5202 0 net490
rlabel metal3 12144 2380 12144 2380 0 net491
rlabel metal1 5336 13974 5336 13974 0 net492
rlabel metal3 17250 12988 17250 12988 0 net493
rlabel metal2 15042 17884 15042 17884 0 net494
rlabel metal1 13156 16014 13156 16014 0 net495
rlabel metal1 15318 11118 15318 11118 0 net496
rlabel metal2 14306 14110 14306 14110 0 net497
rlabel metal1 19734 17204 19734 17204 0 net498
rlabel metal1 25484 10234 25484 10234 0 net499
rlabel metal1 19458 20026 19458 20026 0 net5
rlabel metal1 15916 8398 15916 8398 0 net50
rlabel metal1 6440 12206 6440 12206 0 net500
rlabel metal1 6716 14586 6716 14586 0 net501
rlabel metal1 23460 37230 23460 37230 0 net502
rlabel metal1 22586 37094 22586 37094 0 net503
rlabel metal1 9200 4114 9200 4114 0 net504
rlabel metal1 10442 5746 10442 5746 0 net505
rlabel metal2 12650 20026 12650 20026 0 net506
rlabel metal1 19826 13226 19826 13226 0 net507
rlabel metal2 25254 14620 25254 14620 0 net508
rlabel via1 22034 26299 22034 26299 0 net509
rlabel metal1 20976 14246 20976 14246 0 net51
rlabel metal2 5382 12172 5382 12172 0 net510
rlabel metal1 11822 37978 11822 37978 0 net511
rlabel metal1 13340 21998 13340 21998 0 net512
rlabel metal2 8878 10914 8878 10914 0 net513
rlabel metal2 15318 18054 15318 18054 0 net514
rlabel metal1 11638 24582 11638 24582 0 net515
rlabel metal2 21482 17408 21482 17408 0 net516
rlabel metal1 12006 26962 12006 26962 0 net517
rlabel metal1 16560 29138 16560 29138 0 net518
rlabel metal4 12788 14824 12788 14824 0 net519
rlabel metal1 15318 8874 15318 8874 0 net52
rlabel metal1 17756 20910 17756 20910 0 net520
rlabel metal1 8510 10234 8510 10234 0 net521
rlabel metal1 14674 20944 14674 20944 0 net522
rlabel metal2 6302 13702 6302 13702 0 net523
rlabel metal2 7498 25228 7498 25228 0 net524
rlabel metal1 9982 26554 9982 26554 0 net525
rlabel metal1 8556 23290 8556 23290 0 net526
rlabel metal2 11270 31110 11270 31110 0 net527
rlabel metal1 9108 14518 9108 14518 0 net528
rlabel metal1 17526 18734 17526 18734 0 net529
rlabel metal2 2438 2958 2438 2958 0 net53
rlabel metal1 12282 31348 12282 31348 0 net530
rlabel metal1 17112 13294 17112 13294 0 net531
rlabel metal1 7130 4114 7130 4114 0 net532
rlabel metal2 6026 19958 6026 19958 0 net533
rlabel metal1 18308 38318 18308 38318 0 net534
rlabel metal1 5658 19856 5658 19856 0 net535
rlabel metal2 13570 9146 13570 9146 0 net536
rlabel metal1 15594 18326 15594 18326 0 net537
rlabel metal1 5750 20944 5750 20944 0 net538
rlabel metal2 6946 15436 6946 15436 0 net539
rlabel metal1 18308 9554 18308 9554 0 net54
rlabel metal1 7728 17646 7728 17646 0 net540
rlabel metal2 6762 13770 6762 13770 0 net541
rlabel metal1 8556 4794 8556 4794 0 net542
rlabel metal1 6256 2414 6256 2414 0 net543
rlabel metal1 1610 5168 1610 5168 0 net544
rlabel metal2 4048 4692 4048 4692 0 net545
rlabel metal1 2070 7514 2070 7514 0 net546
rlabel metal1 3726 5882 3726 5882 0 net547
rlabel metal2 24702 52666 24702 52666 0 net548
rlabel metal1 24288 53074 24288 53074 0 net549
rlabel metal1 10028 18326 10028 18326 0 net55
rlabel metal2 24610 53754 24610 53754 0 net550
rlabel metal1 23414 52462 23414 52462 0 net551
rlabel metal1 23368 51986 23368 51986 0 net552
rlabel metal2 2714 3179 2714 3179 0 net56
rlabel metal1 2898 2380 2898 2380 0 net57
rlabel metal2 21298 1768 21298 1768 0 net58
rlabel metal3 5612 12444 5612 12444 0 net59
rlabel via2 15778 17867 15778 17867 0 net6
rlabel metal1 1886 11832 1886 11832 0 net60
rlabel metal2 12650 4896 12650 4896 0 net61
rlabel via2 5474 2499 5474 2499 0 net62
rlabel metal1 12880 46478 12880 46478 0 net63
rlabel metal1 14628 47090 14628 47090 0 net64
rlabel metal2 15686 50218 15686 50218 0 net65
rlabel metal2 17158 49912 17158 49912 0 net66
rlabel metal1 18170 54128 18170 54128 0 net67
rlabel metal3 20447 1156 20447 1156 0 net68
rlabel metal2 24610 50592 24610 50592 0 net69
rlabel metal1 25438 39338 25438 39338 0 net7
rlabel metal1 22080 44166 22080 44166 0 net70
rlabel metal1 21988 51918 21988 51918 0 net71
rlabel metal1 20838 51850 20838 51850 0 net72
rlabel metal1 19090 54026 19090 54026 0 net73
rlabel metal1 21022 52938 21022 52938 0 net74
rlabel metal1 20470 49402 20470 49402 0 net75
rlabel metal1 20332 41446 20332 41446 0 net76
rlabel metal1 18446 8432 18446 8432 0 net77
rlabel metal2 5566 52088 5566 52088 0 net78
rlabel metal2 17526 7905 17526 7905 0 net79
rlabel metal3 16767 35836 16767 35836 0 net8
rlabel via2 13386 13685 13386 13685 0 net80
rlabel metal1 1794 9486 1794 9486 0 net81
rlabel via2 3634 10557 3634 10557 0 net82
rlabel metal2 21022 12087 21022 12087 0 net83
rlabel metal3 13524 14008 13524 14008 0 net84
rlabel metal1 18262 14042 18262 14042 0 net85
rlabel metal1 20930 16762 20930 16762 0 net86
rlabel metal1 16422 15640 16422 15640 0 net87
rlabel metal1 19274 16524 19274 16524 0 net88
rlabel metal2 23966 15062 23966 15062 0 net89
rlabel metal1 25668 40358 25668 40358 0 net9
rlabel metal2 9798 2006 9798 2006 0 net90
rlabel metal1 22402 13498 22402 13498 0 net91
rlabel via2 4738 18173 4738 18173 0 net92
rlabel metal2 20838 19873 20838 19873 0 net93
rlabel metal2 22218 19244 22218 19244 0 net94
rlabel metal1 20884 18938 20884 18938 0 net95
rlabel metal2 23782 21386 23782 21386 0 net96
rlabel metal2 6302 23137 6302 23137 0 net97
rlabel metal2 21850 22066 21850 22066 0 net98
rlabel metal2 21758 26384 21758 26384 0 net99
rlabel metal1 18216 24106 18216 24106 0 prog_clk
rlabel metal2 24242 493 24242 493 0 prog_reset
rlabel metal2 24978 50711 24978 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 24978 51323 24978 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24978 52105 24978 52105 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 24610 52275 24610 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 22678 54026 22678 54026 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 22862 53873 22862 53873 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 24388 55420 24388 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 25262 56236 25262 56236 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 20378 54648 20378 54648 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21758 55711 21758 55711 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 22954 56236 22954 56236 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 24518 53288 24518 53288 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 2683 1836 2683 1836 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 19044 46478 19044 46478 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 25622 33626 25622 33626 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 25024 33490 25024 33490 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 17940 11662 17940 11662 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal1 21022 19142 21022 19142 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal1 20516 15878 20516 15878 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal2 21574 18394 21574 18394 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal1 24978 15470 24978 15470 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal2 6486 24004 6486 24004 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 20838 20468 20838 20468 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 24196 26418 24196 26418 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 21298 24174 21298 24174 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal1 24104 18802 24104 18802 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal2 19090 25738 19090 25738 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal2 21206 27540 21206 27540 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal2 18906 27642 18906 27642 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal2 19366 28866 19366 28866 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal2 18814 32402 18814 32402 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 19596 30702 19596 30702 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 2116 8534 2116 8534 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal2 17020 14348 17020 14348 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 21022 31994 21022 31994 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal2 22586 32028 22586 32028 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 23966 27506 23966 27506 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 23000 34578 23000 34578 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 24932 38930 24932 38930 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 24748 36754 24748 36754 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 23874 37842 23874 37842 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal2 23322 34102 23322 34102 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 20654 33626 20654 33626 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal2 23414 34238 23414 34238 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 21298 33014 21298 33014 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 21206 34850 21206 34850 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal1 24656 19278 24656 19278 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 8602 21386 8602 21386 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 22080 17646 22080 17646 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 19918 23630 19918 23630 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal2 21252 20740 21252 20740 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 18538 21998 18538 21998 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 11684 25874 11684 25874 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal1 21482 43622 21482 43622 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal2 14214 19210 14214 19210 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal1 10534 24582 10534 24582 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 9292 18802 9292 18802 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal2 9614 24548 9614 24548 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 9108 22406 9108 22406 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal1 12627 19278 12627 19278 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 9062 19448 9062 19448 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 15640 21522 15640 21522 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal2 13386 19533 13386 19533 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal2 14674 20604 14674 20604 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 14628 17102 14628 17102 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal1 13110 15878 13110 15878 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 13708 18598 13708 18598 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal2 11178 27948 11178 27948 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal1 12788 28730 12788 28730 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal1 10396 25466 10396 25466 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 9798 9350 9798 9350 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal2 11178 12517 11178 12517 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 6946 7446 6946 7446 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal1 10580 8330 10580 8330 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal1 12328 6834 12328 6834 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 9982 6426 9982 6426 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 15778 13804 15778 13804 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal1 15318 11730 15318 11730 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 16376 19346 16376 19346 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 14674 17680 14674 17680 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal1 18538 19890 18538 19890 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 16100 20230 16100 20230 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal2 18630 16354 18630 16354 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 17618 14926 17618 14926 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal1 15962 9894 15962 9894 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 12834 7378 12834 7378 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal2 14858 4828 14858 4828 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 14582 6222 14582 6222 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16514 4658 16514 4658 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15778 3706 15778 3706 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 14582 28186 14582 28186 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal2 16514 30498 16514 30498 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 13478 31790 13478 31790 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal2 19642 7072 19642 7072 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal2 17802 5406 17802 5406 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal1 21298 10540 21298 10540 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal1 11546 1122 11546 1122 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 20056 13838 20056 13838 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal2 20378 18717 20378 18717 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal2 21666 14841 21666 14841 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 20700 22066 20700 22066 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20976 13362 20976 13362 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal2 16330 21148 16330 21148 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal1 18952 19754 18952 19754 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal2 21482 12665 21482 12665 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal2 18814 22729 18814 22729 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal2 9246 7548 9246 7548 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal1 16652 4046 16652 4046 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal2 17802 4199 17802 4199 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 17112 6222 17112 6222 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal2 20010 4505 20010 4505 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 17802 8806 17802 8806 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal1 13524 23154 13524 23154 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal1 17066 28594 17066 28594 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal2 11730 25228 11730 25228 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal1 15686 26894 15686 26894 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal1 11178 25704 11178 25704 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal1 2208 5678 2208 5678 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20792 18598 20792 18598 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20102 18734 20102 18734 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20194 18326 20194 18326 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 1564 6766 1564 6766 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 24840 26486 24840 26486 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6578 16218 6578 16218 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel via3 1725 4012 1725 4012 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 23368 23834 23368 23834 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15134 22831 15134 22831 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16836 7990 16836 7990 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal2 23414 23307 23414 23307 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19964 17238 19964 17238 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9108 15674 9108 15674 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 21022 24616 21022 24616 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 18538 24667 18538 24667 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4968 6358 4968 6358 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 19596 26010 19596 26010 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 18078 25755 18078 25755 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14490 4488 14490 4488 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 18952 28526 18952 28526 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13478 28560 13478 28560 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14168 6698 14168 6698 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal2 25070 19159 25070 19159 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4462 14790 4462 14790 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3036 8534 3036 8534 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal1 21390 31858 21390 31858 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 17779 13668 17779 13668 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8924 15300 8924 15300 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal2 23920 31756 23920 31756 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 5520 23460 5520 23460 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15134 17204 15134 17204 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 24656 28050 24656 28050 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10994 27421 10994 27421 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal4 14996 19312 14996 19312 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal2 22494 30787 22494 30787 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 22034 29019 22034 29019 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13570 19788 13570 19788 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal1 21528 35462 21528 35462 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18952 29750 18952 29750 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 16031 20876 16031 20876 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 20332 29614 20332 29614 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 21590 19458 21590 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19366 8806 19366 8806 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 24656 22950 24656 22950 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal4 20608 14620 20608 14620 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 2482 17526 2482 0 sb_0__8_.mux_bottom_track_51.out
rlabel via2 22954 17323 22954 17323 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 22494 17051 22494 17051 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2162 9214 2162 9214 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal1 20470 22746 20470 22746 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 22746 19688 22746 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19550 20026 19550 20026 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 2047 8364 2047 8364 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22448 20570 22448 20570 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 22034 20315 22034 20315 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13570 25840 13570 25840 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 15088 32742 15088 32742 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15640 28390 15640 28390 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13064 26350 13064 26350 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10304 26282 10304 26282 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 13478 25874 13478 25874 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 21206 18734 21206 18734 0 sb_0__8_.mux_right_track_10.out
rlabel metal2 13386 23630 13386 23630 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12236 22746 12236 22746 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11408 22406 11408 22406 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7452 12614 7452 12614 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13294 20366 13294 20366 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18722 18734 18722 18734 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 12834 19346 12834 19346 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12650 19380 12650 19380 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15226 19108 15226 19108 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 3726 20570 3726 20570 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 16514 21998 16514 21998 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 18360 12926 18360 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15962 21896 15962 21896 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 4554 18462 4554 18462 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 16330 19754 16330 19754 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14720 17306 14720 17306 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13938 19312 13938 19312 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21942 15623 21942 15623 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 13892 15402 13892 15402 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8234 16728 8234 16728 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16146 26792 16146 26792 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 15180 29478 15180 29478 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15870 28492 15870 28492 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13478 27744 13478 27744 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11822 27030 11822 27030 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16330 27030 16330 27030 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 20792 13906 20792 13906 0 sb_0__8_.mux_right_track_20.out
rlabel metal1 11546 9962 11546 9962 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12190 8772 12190 8772 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16698 16269 16698 16269 0 sb_0__8_.mux_right_track_22.out
rlabel metal2 12834 6766 12834 6766 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12098 7718 12098 7718 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7084 14484 7084 14484 0 sb_0__8_.mux_right_track_24.out
rlabel metal1 11868 6086 11868 6086 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 14306 7701 14306 7701 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2346 13906 2346 13906 0 sb_0__8_.mux_right_track_26.out
rlabel metal1 14536 12614 14536 12614 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 13923 15226 13923 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3956 16150 3956 16150 0 sb_0__8_.mux_right_track_28.out
rlabel metal2 16514 20876 16514 20876 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14352 15130 14352 15130 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16054 18360 16054 18360 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 2668 14382 2668 14382 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 18308 19822 18308 19822 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 15318 15963 15318 15963 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17618 19737 17618 19737 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 3634 13294 3634 13294 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 18630 17646 18630 17646 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 15130 17618 15130 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17894 17357 17894 17357 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4094 10710 4094 10710 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 16652 11118 16652 11118 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16422 11152 16422 11152 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4922 11186 4922 11186 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9108 4794 9108 4794 0 sb_0__8_.mux_right_track_36.out
rlabel metal2 15962 5746 15962 5746 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15502 4896 15502 4896 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 1610 11016 1610 11016 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 15548 6426 15548 6426 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1748 12682 1748 12682 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 21574 20876 21574 20876 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 15502 27302 15502 27302 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15272 27438 15272 27438 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 25330 14904 25330 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14536 25194 14536 25194 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21482 24480 21482 24480 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 4462 8534 4462 8534 0 sb_0__8_.mux_right_track_40.out
rlabel metal1 20240 6222 20240 6222 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20516 6086 20516 6086 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1978 12104 1978 12104 0 sb_0__8_.mux_right_track_42.out
rlabel metal1 19688 10778 19688 10778 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 2162 12189 2162 12189 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 3818 10302 3818 10302 0 sb_0__8_.mux_right_track_44.out
rlabel metal1 19826 14042 19826 14042 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19550 13906 19550 13906 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14214 12784 14214 12784 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4646 9622 4646 9622 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 20332 21862 20332 21862 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20286 13498 20286 13498 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16238 15810 16238 15810 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 4738 8500 4738 8500 0 sb_0__8_.mux_right_track_48.out
rlabel metal2 21206 15130 21206 15130 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 11322 20378 11322 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2714 9401 2714 9401 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 17204 884 17204 884 0 sb_0__8_.mux_right_track_50.out
rlabel metal2 22586 13872 22586 13872 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20700 4046 20700 4046 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6348 4250 6348 4250 0 sb_0__8_.mux_right_track_52.out
rlabel metal1 24564 5746 24564 5746 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24610 5593 24610 5593 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8280 3706 8280 3706 0 sb_0__8_.mux_right_track_54.out
rlabel metal1 17894 4114 17894 4114 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16790 3774 16790 3774 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6348 2618 6348 2618 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 17572 6426 17572 6426 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9338 1938 9338 1938 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9706 8602 9706 8602 0 sb_0__8_.mux_right_track_58.out
rlabel metal1 17250 16966 17250 16966 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 11220 13202 11220 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16882 11832 16882 11832 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7682 23460 7682 23460 0 sb_0__8_.mux_right_track_6.out
rlabel metal1 16100 26010 16100 26010 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15410 25840 15410 25840 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14122 22950 14122 22950 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 22984 12742 22984 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12006 23664 12006 23664 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18676 19482 18676 19482 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 13294 25075 13294 25075 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13202 24956 13202 24956 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 23834 12558 23834 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10028 23154 10028 23154 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11730 22984 11730 22984 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
