magic
tech sky130A
magscale 1 2
timestamp 1680088070
<< viali >>
rect 3985 24361 4019 24395
rect 11713 24361 11747 24395
rect 14289 24361 14323 24395
rect 38577 24361 38611 24395
rect 42165 24361 42199 24395
rect 44741 24361 44775 24395
rect 29009 24293 29043 24327
rect 31309 24293 31343 24327
rect 32781 24293 32815 24327
rect 33517 24293 33551 24327
rect 36829 24293 36863 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 16865 24225 16899 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25145 24225 25179 24259
rect 26341 24225 26375 24259
rect 27721 24225 27755 24259
rect 29745 24225 29779 24259
rect 34253 24225 34287 24259
rect 37013 24225 37047 24259
rect 40049 24225 40083 24259
rect 40325 24225 40359 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 15117 24157 15151 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22017 24157 22051 24191
rect 24041 24157 24075 24191
rect 27629 24157 27663 24191
rect 28549 24157 28583 24191
rect 29193 24157 29227 24191
rect 30021 24157 30055 24191
rect 31493 24157 31527 24191
rect 32505 24157 32539 24191
rect 33333 24157 33367 24191
rect 34069 24157 34103 24191
rect 34989 24157 35023 24191
rect 35725 24157 35759 24191
rect 36553 24157 36587 24191
rect 37657 24157 37691 24191
rect 38485 24157 38519 24191
rect 39221 24157 39255 24191
rect 41521 24157 41555 24191
rect 41797 24157 41831 24191
rect 42625 24157 42659 24191
rect 45201 24157 45235 24191
rect 45937 24157 45971 24191
rect 46673 24157 46707 24191
rect 47225 24157 47259 24191
rect 47777 24157 47811 24191
rect 48513 24157 48547 24191
rect 49065 24157 49099 24191
rect 17141 24089 17175 24123
rect 18981 24089 19015 24123
rect 26249 24089 26283 24123
rect 35909 24089 35943 24123
rect 37933 24089 37967 24123
rect 6561 24021 6595 24055
rect 9137 24021 9171 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 23857 24021 23891 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 25053 24021 25087 24055
rect 25789 24021 25823 24055
rect 26157 24021 26191 24055
rect 27169 24021 27203 24055
rect 27537 24021 27571 24055
rect 28365 24021 28399 24055
rect 30849 24021 30883 24055
rect 31769 24021 31803 24055
rect 32321 24021 32355 24055
rect 35081 24021 35115 24055
rect 36369 24021 36403 24055
rect 37473 24021 37507 24055
rect 39313 24021 39347 24055
rect 41337 24021 41371 24055
rect 43913 24021 43947 24055
rect 45385 24021 45419 24055
rect 46121 24021 46155 24055
rect 46857 24021 46891 24055
rect 47961 24021 47995 24055
rect 48697 24021 48731 24055
rect 49525 24021 49559 24055
rect 12357 23817 12391 23851
rect 21097 23817 21131 23851
rect 24225 23817 24259 23851
rect 30941 23817 30975 23851
rect 31309 23817 31343 23851
rect 32965 23817 32999 23851
rect 34069 23817 34103 23851
rect 34805 23817 34839 23851
rect 38485 23817 38519 23851
rect 39037 23817 39071 23851
rect 39865 23817 39899 23851
rect 43269 23817 43303 23851
rect 45753 23817 45787 23851
rect 47593 23817 47627 23851
rect 3985 23749 4019 23783
rect 7205 23749 7239 23783
rect 9137 23749 9171 23783
rect 10977 23749 11011 23783
rect 14197 23749 14231 23783
rect 16129 23749 16163 23783
rect 18981 23749 19015 23783
rect 21557 23749 21591 23783
rect 30113 23749 30147 23783
rect 33425 23749 33459 23783
rect 35449 23749 35483 23783
rect 35633 23749 35667 23783
rect 2145 23681 2179 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 7113 23681 7147 23715
rect 8125 23681 8159 23715
rect 9873 23681 9907 23715
rect 11805 23681 11839 23715
rect 12265 23681 12299 23715
rect 13093 23681 13127 23715
rect 14933 23681 14967 23715
rect 17049 23681 17083 23715
rect 18705 23681 18739 23715
rect 21005 23681 21039 23715
rect 29561 23681 29595 23715
rect 31493 23681 31527 23715
rect 33977 23681 34011 23715
rect 34713 23681 34747 23715
rect 36277 23681 36311 23715
rect 36921 23681 36955 23715
rect 37289 23681 37323 23715
rect 37933 23681 37967 23715
rect 38209 23681 38243 23715
rect 41521 23681 41555 23715
rect 41797 23681 41831 23715
rect 43545 23681 43579 23715
rect 44281 23681 44315 23715
rect 44833 23681 44867 23715
rect 46765 23681 46799 23715
rect 47317 23681 47351 23715
rect 48053 23681 48087 23715
rect 48329 23681 48363 23715
rect 49065 23681 49099 23715
rect 5457 23613 5491 23647
rect 7389 23613 7423 23647
rect 12541 23613 12575 23647
rect 17877 23613 17911 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 30665 23613 30699 23647
rect 32321 23613 32355 23647
rect 6561 23545 6595 23579
rect 23765 23545 23799 23579
rect 29377 23545 29411 23579
rect 31769 23545 31803 23579
rect 32137 23545 32171 23579
rect 37749 23545 37783 23579
rect 41337 23545 41371 23579
rect 2237 23477 2271 23511
rect 6377 23477 6411 23511
rect 6745 23477 6779 23511
rect 11529 23477 11563 23511
rect 11897 23477 11931 23511
rect 20453 23477 20487 23511
rect 26617 23477 26651 23511
rect 28917 23477 28951 23511
rect 30205 23477 30239 23511
rect 30757 23477 30791 23511
rect 36093 23477 36127 23511
rect 36737 23477 36771 23511
rect 43729 23477 43763 23511
rect 44465 23477 44499 23511
rect 46949 23477 46983 23511
rect 48513 23477 48547 23511
rect 49249 23477 49283 23511
rect 14473 23273 14507 23307
rect 27524 23273 27558 23307
rect 29009 23273 29043 23307
rect 30002 23273 30036 23307
rect 31953 23273 31987 23307
rect 32505 23273 32539 23307
rect 36645 23273 36679 23307
rect 36829 23273 36863 23307
rect 37289 23273 37323 23307
rect 4169 23205 4203 23239
rect 18889 23205 18923 23239
rect 25789 23205 25823 23239
rect 34345 23205 34379 23239
rect 36001 23205 36035 23239
rect 4813 23137 4847 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11529 23137 11563 23171
rect 16497 23137 16531 23171
rect 20085 23137 20119 23171
rect 21833 23137 21867 23171
rect 22569 23137 22603 23171
rect 25145 23137 25179 23171
rect 26341 23137 26375 23171
rect 27261 23137 27295 23171
rect 29377 23137 29411 23171
rect 29745 23137 29779 23171
rect 1777 23069 1811 23103
rect 3617 23069 3651 23103
rect 4629 23069 4663 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 19625 23069 19659 23103
rect 22293 23069 22327 23103
rect 33333 23069 33367 23103
rect 34069 23069 34103 23103
rect 35081 23069 35115 23103
rect 35725 23069 35759 23103
rect 36185 23069 36219 23103
rect 48605 23069 48639 23103
rect 49065 23069 49099 23103
rect 2789 23001 2823 23035
rect 9597 23001 9631 23035
rect 11805 23001 11839 23035
rect 13645 23001 13679 23035
rect 13829 23001 13863 23035
rect 14381 23001 14415 23035
rect 17417 23001 17451 23035
rect 20361 23001 20395 23035
rect 26249 23001 26283 23035
rect 32413 23001 32447 23035
rect 33149 23001 33183 23035
rect 33885 23001 33919 23035
rect 3801 22933 3835 22967
rect 4077 22933 4111 22967
rect 4537 22933 4571 22967
rect 9045 22933 9079 22967
rect 11069 22933 11103 22967
rect 13277 22933 13311 22967
rect 14933 22933 14967 22967
rect 19441 22933 19475 22967
rect 24041 22933 24075 22967
rect 24593 22933 24627 22967
rect 24961 22933 24995 22967
rect 25053 22933 25087 22967
rect 26157 22933 26191 22967
rect 26801 22933 26835 22967
rect 31493 22933 31527 22967
rect 31769 22933 31803 22967
rect 34897 22933 34931 22967
rect 35541 22933 35575 22967
rect 48421 22933 48455 22967
rect 49249 22933 49283 22967
rect 14657 22729 14691 22763
rect 21465 22729 21499 22763
rect 22477 22729 22511 22763
rect 25789 22729 25823 22763
rect 32505 22729 32539 22763
rect 33149 22729 33183 22763
rect 39957 22729 39991 22763
rect 48697 22729 48731 22763
rect 49341 22729 49375 22763
rect 10701 22661 10735 22695
rect 11805 22661 11839 22695
rect 16129 22661 16163 22695
rect 17141 22661 17175 22695
rect 23397 22661 23431 22695
rect 28641 22661 28675 22695
rect 31033 22661 31067 22695
rect 1777 22593 1811 22627
rect 3801 22593 3835 22627
rect 4813 22593 4847 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 7941 22593 7975 22627
rect 9965 22593 9999 22627
rect 15117 22593 15151 22627
rect 19257 22593 19291 22627
rect 19717 22593 19751 22627
rect 23121 22593 23155 22627
rect 25697 22593 25731 22627
rect 26341 22593 26375 22627
rect 27537 22593 27571 22627
rect 30941 22593 30975 22627
rect 31769 22593 31803 22627
rect 32413 22593 32447 22627
rect 33609 22593 33643 22627
rect 33885 22593 33919 22627
rect 37841 22593 37875 22627
rect 2789 22525 2823 22559
rect 3893 22525 3927 22559
rect 4077 22525 4111 22559
rect 5089 22525 5123 22559
rect 7389 22525 7423 22559
rect 8677 22525 8711 22559
rect 12449 22525 12483 22559
rect 12725 22525 12759 22559
rect 16865 22525 16899 22559
rect 19993 22525 20027 22559
rect 24869 22525 24903 22559
rect 25881 22525 25915 22559
rect 27629 22525 27663 22559
rect 27721 22525 27755 22559
rect 28365 22525 28399 22559
rect 31125 22525 31159 22559
rect 31585 22525 31619 22559
rect 38117 22525 38151 22559
rect 18613 22457 18647 22491
rect 27169 22457 27203 22491
rect 35357 22457 35391 22491
rect 3433 22389 3467 22423
rect 6377 22389 6411 22423
rect 6745 22389 6779 22423
rect 11897 22389 11931 22423
rect 14197 22389 14231 22423
rect 19073 22389 19107 22423
rect 22017 22389 22051 22423
rect 22109 22389 22143 22423
rect 25329 22389 25363 22423
rect 26525 22389 26559 22423
rect 26709 22389 26743 22423
rect 30113 22389 30147 22423
rect 30573 22389 30607 22423
rect 32873 22389 32907 22423
rect 33333 22389 33367 22423
rect 34713 22389 34747 22423
rect 34897 22389 34931 22423
rect 39589 22389 39623 22423
rect 49525 22389 49559 22423
rect 18889 22185 18923 22219
rect 22201 22185 22235 22219
rect 10241 22117 10275 22151
rect 27537 22117 27571 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 9229 22049 9263 22083
rect 9965 22049 9999 22083
rect 11253 22049 11287 22083
rect 13369 22049 13403 22083
rect 14565 22049 14599 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 20913 22049 20947 22083
rect 23949 22049 23983 22083
rect 25145 22049 25179 22083
rect 26065 22049 26099 22083
rect 27997 22049 28031 22083
rect 30757 22049 30791 22083
rect 31585 22049 31619 22083
rect 33701 22049 33735 22083
rect 1777 21981 1811 22015
rect 4077 21981 4111 22015
rect 6285 21981 6319 22015
rect 7021 21981 7055 22015
rect 8769 21981 8803 22015
rect 10701 21981 10735 22015
rect 12541 21981 12575 22015
rect 14381 21981 14415 22015
rect 15393 21981 15427 22015
rect 20361 21981 20395 22015
rect 23765 21981 23799 22015
rect 25789 21981 25823 22015
rect 28825 21981 28859 22015
rect 29285 21981 29319 22015
rect 29837 21981 29871 22015
rect 30573 21981 30607 22015
rect 32597 21981 32631 22015
rect 32873 21981 32907 22015
rect 49065 21981 49099 22015
rect 3617 21913 3651 21947
rect 7849 21913 7883 21947
rect 8585 21913 8619 21947
rect 17417 21913 17451 21947
rect 19533 21913 19567 21947
rect 19993 21913 20027 21947
rect 22661 21913 22695 21947
rect 24961 21913 24995 21947
rect 30481 21913 30515 21947
rect 31401 21913 31435 21947
rect 31861 21913 31895 21947
rect 3341 21845 3375 21879
rect 5825 21845 5859 21879
rect 6101 21845 6135 21879
rect 8953 21845 8987 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 9781 21845 9815 21879
rect 14933 21845 14967 21879
rect 19625 21845 19659 21879
rect 22109 21845 22143 21879
rect 23305 21845 23339 21879
rect 23673 21845 23707 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 28641 21845 28675 21879
rect 29193 21845 29227 21879
rect 29561 21845 29595 21879
rect 30113 21845 30147 21879
rect 32137 21845 32171 21879
rect 49249 21845 49283 21879
rect 9413 21641 9447 21675
rect 9873 21641 9907 21675
rect 15485 21641 15519 21675
rect 15945 21641 15979 21675
rect 16037 21641 16071 21675
rect 22477 21641 22511 21675
rect 25973 21641 26007 21675
rect 27261 21641 27295 21675
rect 27721 21641 27755 21675
rect 4353 21573 4387 21607
rect 7021 21573 7055 21607
rect 7941 21573 7975 21607
rect 13369 21573 13403 21607
rect 23673 21573 23707 21607
rect 26065 21573 26099 21607
rect 31125 21573 31159 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 5641 21505 5675 21539
rect 10241 21505 10275 21539
rect 10701 21505 10735 21539
rect 11161 21505 11195 21539
rect 11253 21505 11287 21539
rect 12173 21505 12207 21539
rect 13093 21505 13127 21539
rect 17049 21505 17083 21539
rect 21281 21505 21315 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 26709 21505 26743 21539
rect 27629 21505 27663 21539
rect 28457 21505 28491 21539
rect 31033 21505 31067 21539
rect 31769 21505 31803 21539
rect 32413 21505 32447 21539
rect 47961 21505 47995 21539
rect 2053 21437 2087 21471
rect 5733 21437 5767 21471
rect 5917 21437 5951 21471
rect 7654 21437 7688 21471
rect 10333 21437 10367 21471
rect 10425 21437 10459 21471
rect 10977 21437 11011 21471
rect 12265 21437 12299 21471
rect 12357 21437 12391 21471
rect 16221 21437 16255 21471
rect 17325 21437 17359 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 22661 21437 22695 21471
rect 25145 21437 25179 21471
rect 26249 21437 26283 21471
rect 27905 21437 27939 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 49157 21437 49191 21471
rect 7205 21369 7239 21403
rect 15209 21369 15243 21403
rect 15577 21369 15611 21403
rect 22017 21369 22051 21403
rect 5273 21301 5307 21335
rect 6377 21301 6411 21335
rect 6653 21301 6687 21335
rect 9781 21301 9815 21335
rect 11805 21301 11839 21335
rect 14841 21301 14875 21335
rect 20453 21301 20487 21335
rect 20729 21301 20763 21335
rect 21005 21301 21039 21335
rect 23029 21301 23063 21335
rect 25605 21301 25639 21335
rect 30205 21301 30239 21335
rect 30665 21301 30699 21335
rect 31861 21301 31895 21335
rect 32505 21301 32539 21335
rect 47685 21301 47719 21335
rect 13829 21097 13863 21131
rect 32505 21097 32539 21131
rect 21649 21029 21683 21063
rect 21833 21029 21867 21063
rect 3893 20961 3927 20995
rect 3985 20961 4019 20995
rect 4261 20961 4295 20995
rect 5733 20961 5767 20995
rect 8493 20961 8527 20995
rect 12541 20961 12575 20995
rect 13737 20961 13771 20995
rect 14197 20961 14231 20995
rect 15117 20961 15151 20995
rect 16405 20961 16439 20995
rect 17601 20961 17635 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 19717 20961 19751 20995
rect 22753 20961 22787 20995
rect 23857 20961 23891 20995
rect 25145 20961 25179 20995
rect 25329 20961 25363 20995
rect 26065 20961 26099 20995
rect 28549 20961 28583 20995
rect 30021 20961 30055 20995
rect 1777 20893 1811 20927
rect 5457 20893 5491 20927
rect 9321 20893 9355 20927
rect 10977 20893 11011 20927
rect 12081 20893 12115 20927
rect 15025 20893 15059 20927
rect 16221 20893 16255 20927
rect 17417 20893 17451 20927
rect 18521 20893 18555 20927
rect 19441 20893 19475 20927
rect 28273 20893 28307 20927
rect 29745 20893 29779 20927
rect 31861 20893 31895 20927
rect 32689 20893 32723 20927
rect 2789 20825 2823 20859
rect 8217 20825 8251 20859
rect 10057 20825 10091 20859
rect 11345 20825 11379 20859
rect 22477 20825 22511 20859
rect 23673 20825 23707 20859
rect 25053 20825 25087 20859
rect 26341 20825 26375 20859
rect 31125 20825 31159 20859
rect 5181 20757 5215 20791
rect 7205 20757 7239 20791
rect 7481 20757 7515 20791
rect 7849 20757 7883 20791
rect 8309 20757 8343 20791
rect 11437 20757 11471 20791
rect 14565 20757 14599 20791
rect 14933 20757 14967 20791
rect 15761 20757 15795 20791
rect 16129 20757 16163 20791
rect 16957 20757 16991 20791
rect 17325 20757 17359 20791
rect 18153 20757 18187 20791
rect 21189 20757 21223 20791
rect 22109 20757 22143 20791
rect 22569 20757 22603 20791
rect 23305 20757 23339 20791
rect 23765 20757 23799 20791
rect 24685 20757 24719 20791
rect 25789 20757 25823 20791
rect 27813 20757 27847 20791
rect 31217 20757 31251 20791
rect 31953 20757 31987 20791
rect 13001 20553 13035 20587
rect 16129 20553 16163 20587
rect 17509 20553 17543 20587
rect 18521 20553 18555 20587
rect 18889 20553 18923 20587
rect 18981 20553 19015 20587
rect 23397 20553 23431 20587
rect 27537 20553 27571 20587
rect 27629 20553 27663 20587
rect 31033 20553 31067 20587
rect 8769 20485 8803 20519
rect 22017 20485 22051 20519
rect 22753 20485 22787 20519
rect 28641 20485 28675 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5641 20417 5675 20451
rect 6561 20417 6595 20451
rect 8401 20417 8435 20451
rect 11805 20417 11839 20451
rect 12909 20417 12943 20451
rect 13461 20417 13495 20451
rect 13737 20417 13771 20451
rect 16037 20417 16071 20451
rect 17417 20417 17451 20451
rect 19717 20417 19751 20451
rect 24317 20417 24351 20451
rect 26433 20417 26467 20451
rect 26709 20417 26743 20451
rect 28365 20417 28399 20451
rect 30941 20417 30975 20451
rect 31585 20417 31619 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 5733 20349 5767 20383
rect 5825 20349 5859 20383
rect 7021 20349 7055 20383
rect 9413 20349 9447 20383
rect 9689 20349 9723 20383
rect 11161 20349 11195 20383
rect 12449 20349 12483 20383
rect 13185 20349 13219 20383
rect 14013 20349 14047 20383
rect 16773 20349 16807 20383
rect 17601 20349 17635 20383
rect 19073 20349 19107 20383
rect 19993 20349 20027 20383
rect 24041 20349 24075 20383
rect 24593 20349 24627 20383
rect 26065 20349 26099 20383
rect 27721 20349 27755 20383
rect 31125 20349 31159 20383
rect 8953 20281 8987 20315
rect 5273 20213 5307 20247
rect 11897 20213 11931 20247
rect 12541 20213 12575 20247
rect 13645 20213 13679 20247
rect 15485 20213 15519 20247
rect 17049 20213 17083 20247
rect 18245 20213 18279 20247
rect 21465 20213 21499 20247
rect 27169 20213 27203 20247
rect 30113 20213 30147 20247
rect 30573 20213 30607 20247
rect 10885 20009 10919 20043
rect 11161 20009 11195 20043
rect 11529 20009 11563 20043
rect 13001 20009 13035 20043
rect 17233 20009 17267 20043
rect 18705 20009 18739 20043
rect 30757 20009 30791 20043
rect 16957 19941 16991 19975
rect 24685 19941 24719 19975
rect 27629 19941 27663 19975
rect 29745 19941 29779 19975
rect 30481 19941 30515 19975
rect 4537 19873 4571 19907
rect 4813 19873 4847 19907
rect 6745 19873 6779 19907
rect 7021 19873 7055 19907
rect 9137 19873 9171 19907
rect 12357 19873 12391 19907
rect 13645 19873 13679 19907
rect 14841 19873 14875 19907
rect 17877 19873 17911 19907
rect 20545 19873 20579 19907
rect 23857 19873 23891 19907
rect 25145 19873 25179 19907
rect 25329 19873 25363 19907
rect 28365 19873 28399 19907
rect 28641 19873 28675 19907
rect 31309 19873 31343 19907
rect 1777 19805 1811 19839
rect 12173 19805 12207 19839
rect 12265 19805 12299 19839
rect 14565 19805 14599 19839
rect 17693 19805 17727 19839
rect 18889 19805 18923 19839
rect 20269 19805 20303 19839
rect 22569 19805 22603 19839
rect 25881 19805 25915 19839
rect 29929 19805 29963 19839
rect 31125 19805 31159 19839
rect 31217 19805 31251 19839
rect 2789 19737 2823 19771
rect 9413 19737 9447 19771
rect 13369 19737 13403 19771
rect 13461 19737 13495 19771
rect 19625 19737 19659 19771
rect 23765 19737 23799 19771
rect 26157 19737 26191 19771
rect 6285 19669 6319 19703
rect 8493 19669 8527 19703
rect 11805 19669 11839 19703
rect 13921 19669 13955 19703
rect 14197 19669 14231 19703
rect 14473 19669 14507 19703
rect 16313 19669 16347 19703
rect 16773 19669 16807 19703
rect 17601 19669 17635 19703
rect 18429 19669 18463 19703
rect 19717 19669 19751 19703
rect 22017 19669 22051 19703
rect 22661 19669 22695 19703
rect 23305 19669 23339 19703
rect 23673 19669 23707 19703
rect 25053 19669 25087 19703
rect 27905 19669 27939 19703
rect 30297 19669 30331 19703
rect 5273 19465 5307 19499
rect 5733 19465 5767 19499
rect 10425 19465 10459 19499
rect 10885 19465 10919 19499
rect 14841 19465 14875 19499
rect 18337 19465 18371 19499
rect 19073 19465 19107 19499
rect 21465 19465 21499 19499
rect 22385 19465 22419 19499
rect 23673 19465 23707 19499
rect 26433 19465 26467 19499
rect 30481 19465 30515 19499
rect 4353 19397 4387 19431
rect 5641 19397 5675 19431
rect 7481 19397 7515 19431
rect 9321 19397 9355 19431
rect 10149 19397 10183 19431
rect 14289 19397 14323 19431
rect 22477 19397 22511 19431
rect 23121 19397 23155 19431
rect 28549 19397 28583 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 6561 19329 6595 19363
rect 8585 19329 8619 19363
rect 10333 19329 10367 19363
rect 10793 19329 10827 19363
rect 11713 19329 11747 19363
rect 14749 19329 14783 19363
rect 15669 19329 15703 19363
rect 16497 19329 16531 19363
rect 16773 19329 16807 19363
rect 17417 19329 17451 19363
rect 18245 19329 18279 19363
rect 19257 19329 19291 19363
rect 24041 19329 24075 19363
rect 24133 19329 24167 19363
rect 24961 19329 24995 19363
rect 27261 19329 27295 19363
rect 30665 19329 30699 19363
rect 5917 19261 5951 19295
rect 10977 19261 11011 19295
rect 11989 19261 12023 19295
rect 13461 19261 13495 19295
rect 14933 19261 14967 19295
rect 16957 19261 16991 19295
rect 17141 19261 17175 19295
rect 18429 19261 18463 19295
rect 19717 19261 19751 19295
rect 22661 19261 22695 19295
rect 24317 19261 24351 19295
rect 25789 19261 25823 19295
rect 28273 19261 28307 19295
rect 14381 19193 14415 19227
rect 15853 19193 15887 19227
rect 22017 19193 22051 19227
rect 23305 19193 23339 19227
rect 13737 19125 13771 19159
rect 13921 19125 13955 19159
rect 14013 19125 14047 19159
rect 15209 19125 15243 19159
rect 15393 19125 15427 19159
rect 16037 19125 16071 19159
rect 16221 19125 16255 19159
rect 17233 19125 17267 19159
rect 17601 19125 17635 19159
rect 17693 19125 17727 19159
rect 17877 19125 17911 19159
rect 19980 19125 20014 19159
rect 27997 19125 28031 19159
rect 30021 19125 30055 19159
rect 30941 19125 30975 19159
rect 7100 18921 7134 18955
rect 9413 18921 9447 18955
rect 11069 18921 11103 18955
rect 11621 18921 11655 18955
rect 22937 18921 22971 18955
rect 23397 18921 23431 18955
rect 24041 18921 24075 18955
rect 25145 18921 25179 18955
rect 27169 18921 27203 18955
rect 30757 18921 30791 18955
rect 10517 18853 10551 18887
rect 18153 18853 18187 18887
rect 2053 18785 2087 18819
rect 6837 18785 6871 18819
rect 10057 18785 10091 18819
rect 12265 18785 12299 18819
rect 13553 18785 13587 18819
rect 15025 18785 15059 18819
rect 15209 18785 15243 18819
rect 17509 18785 17543 18819
rect 18705 18785 18739 18819
rect 20361 18785 20395 18819
rect 21189 18785 21223 18819
rect 21465 18785 21499 18819
rect 24593 18785 24627 18819
rect 25421 18785 25455 18819
rect 30205 18785 30239 18819
rect 30297 18785 30331 18819
rect 1777 18717 1811 18751
rect 4629 18717 4663 18751
rect 9781 18717 9815 18751
rect 12817 18717 12851 18751
rect 14197 18717 14231 18751
rect 18521 18717 18555 18751
rect 19625 18717 19659 18751
rect 23581 18717 23615 18751
rect 27629 18717 27663 18751
rect 27905 18717 27939 18751
rect 4905 18649 4939 18683
rect 10977 18649 11011 18683
rect 14565 18649 14599 18683
rect 15492 18649 15526 18683
rect 20913 18649 20947 18683
rect 25697 18649 25731 18683
rect 3617 18581 3651 18615
rect 3985 18581 4019 18615
rect 6377 18581 6411 18615
rect 8585 18581 8619 18615
rect 9137 18581 9171 18615
rect 9873 18581 9907 18615
rect 11989 18581 12023 18615
rect 12081 18581 12115 18615
rect 13829 18581 13863 18615
rect 14657 18581 14691 18615
rect 14933 18581 14967 18615
rect 16957 18581 16991 18615
rect 18613 18581 18647 18615
rect 19349 18581 19383 18615
rect 24225 18581 24259 18615
rect 29745 18581 29779 18615
rect 30113 18581 30147 18615
rect 15025 18377 15059 18411
rect 16497 18377 16531 18411
rect 17325 18377 17359 18411
rect 20729 18377 20763 18411
rect 24869 18377 24903 18411
rect 26801 18377 26835 18411
rect 27169 18377 27203 18411
rect 4445 18309 4479 18343
rect 9781 18309 9815 18343
rect 14473 18309 14507 18343
rect 18153 18309 18187 18343
rect 21097 18309 21131 18343
rect 22569 18309 22603 18343
rect 22845 18309 22879 18343
rect 25329 18309 25363 18343
rect 26065 18309 26099 18343
rect 28365 18309 28399 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 5641 18241 5675 18275
rect 5733 18241 5767 18275
rect 6745 18241 6779 18275
rect 8493 18241 8527 18275
rect 10793 18241 10827 18275
rect 12357 18241 12391 18275
rect 12449 18241 12483 18275
rect 13001 18241 13035 18275
rect 13645 18241 13679 18275
rect 15393 18241 15427 18275
rect 17233 18241 17267 18275
rect 19901 18241 19935 18275
rect 21189 18241 21223 18275
rect 26525 18241 26559 18275
rect 28089 18241 28123 18275
rect 30665 18241 30699 18275
rect 2053 18173 2087 18207
rect 5825 18173 5859 18207
rect 7021 18173 7055 18207
rect 9229 18173 9263 18207
rect 10885 18173 10919 18207
rect 10977 18173 11011 18207
rect 12541 18173 12575 18207
rect 15485 18173 15519 18207
rect 15669 18173 15703 18207
rect 17417 18173 17451 18207
rect 18337 18173 18371 18207
rect 18889 18173 18923 18207
rect 19993 18173 20027 18207
rect 20085 18173 20119 18207
rect 21373 18173 21407 18207
rect 22017 18173 22051 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 30757 18173 30791 18207
rect 30849 18173 30883 18207
rect 31401 18173 31435 18207
rect 9873 18105 9907 18139
rect 13277 18105 13311 18139
rect 19533 18105 19567 18139
rect 30297 18105 30331 18139
rect 5273 18037 5307 18071
rect 10425 18037 10459 18071
rect 11989 18037 12023 18071
rect 16037 18037 16071 18071
rect 16221 18037 16255 18071
rect 16865 18037 16899 18071
rect 29837 18037 29871 18071
rect 31585 18037 31619 18071
rect 3617 17833 3651 17867
rect 3893 17833 3927 17867
rect 6653 17833 6687 17867
rect 7849 17833 7883 17867
rect 10609 17833 10643 17867
rect 11621 17833 11655 17867
rect 13737 17833 13771 17867
rect 14473 17833 14507 17867
rect 19671 17833 19705 17867
rect 21833 17833 21867 17867
rect 4445 17765 4479 17799
rect 20729 17765 20763 17799
rect 26617 17765 26651 17799
rect 29745 17765 29779 17799
rect 7389 17697 7423 17731
rect 8309 17697 8343 17731
rect 8401 17697 8435 17731
rect 9873 17697 9907 17731
rect 11161 17697 11195 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 19441 17697 19475 17731
rect 21281 17697 21315 17731
rect 24869 17697 24903 17731
rect 27077 17697 27111 17731
rect 30205 17697 30239 17731
rect 30297 17697 30331 17731
rect 31493 17697 31527 17731
rect 1777 17629 1811 17663
rect 4905 17629 4939 17663
rect 8217 17629 8251 17663
rect 10977 17629 11011 17663
rect 11989 17629 12023 17663
rect 21189 17629 21223 17663
rect 22293 17629 22327 17663
rect 31309 17629 31343 17663
rect 31401 17629 31435 17663
rect 2513 17561 2547 17595
rect 4261 17561 4295 17595
rect 5181 17561 5215 17595
rect 7205 17561 7239 17595
rect 9137 17561 9171 17595
rect 12265 17561 12299 17595
rect 14381 17561 14415 17595
rect 18337 17561 18371 17595
rect 21097 17561 21131 17595
rect 22569 17561 22603 17595
rect 24409 17561 24443 17595
rect 25145 17561 25179 17595
rect 27353 17561 27387 17595
rect 30113 17561 30147 17595
rect 11069 17493 11103 17527
rect 14841 17493 14875 17527
rect 15025 17493 15059 17527
rect 15393 17493 15427 17527
rect 15945 17493 15979 17527
rect 18061 17493 18095 17527
rect 18705 17493 18739 17527
rect 21925 17493 21959 17527
rect 24041 17493 24075 17527
rect 28825 17493 28859 17527
rect 29193 17493 29227 17527
rect 30941 17493 30975 17527
rect 5273 17289 5307 17323
rect 7297 17289 7331 17323
rect 8033 17289 8067 17323
rect 8493 17289 8527 17323
rect 11253 17289 11287 17323
rect 12541 17289 12575 17323
rect 14197 17289 14231 17323
rect 16129 17289 16163 17323
rect 22017 17289 22051 17323
rect 22385 17289 22419 17323
rect 23673 17289 23707 17323
rect 23765 17289 23799 17323
rect 30941 17289 30975 17323
rect 4629 17221 4663 17255
rect 10977 17221 11011 17255
rect 12909 17221 12943 17255
rect 14749 17221 14783 17255
rect 20177 17221 20211 17255
rect 21097 17221 21131 17255
rect 22477 17221 22511 17255
rect 24961 17221 24995 17255
rect 26801 17221 26835 17255
rect 30573 17221 30607 17255
rect 1777 17153 1811 17187
rect 3617 17153 3651 17187
rect 5641 17153 5675 17187
rect 5733 17153 5767 17187
rect 7205 17153 7239 17187
rect 8401 17153 8435 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 10793 17153 10827 17187
rect 11805 17153 11839 17187
rect 14105 17153 14139 17187
rect 15669 17153 15703 17187
rect 16313 17153 16347 17187
rect 17233 17153 17267 17187
rect 24685 17153 24719 17187
rect 27813 17153 27847 17187
rect 30849 17153 30883 17187
rect 2053 17085 2087 17119
rect 5825 17085 5859 17119
rect 7481 17085 7515 17119
rect 8677 17085 8711 17119
rect 10057 17085 10091 17119
rect 13001 17085 13035 17119
rect 13185 17085 13219 17119
rect 14381 17085 14415 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 18153 17085 18187 17119
rect 18429 17085 18463 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 22569 17085 22603 17119
rect 23857 17085 23891 17119
rect 26433 17085 26467 17119
rect 27169 17085 27203 17119
rect 28089 17085 28123 17119
rect 6837 17017 6871 17051
rect 13737 17017 13771 17051
rect 16865 17017 16899 17051
rect 20729 17017 20763 17051
rect 6561 16949 6595 16983
rect 9045 16949 9079 16983
rect 9505 16949 9539 16983
rect 11897 16949 11931 16983
rect 15485 16949 15519 16983
rect 19901 16949 19935 16983
rect 20361 16949 20395 16983
rect 23305 16949 23339 16983
rect 24409 16949 24443 16983
rect 29561 16949 29595 16983
rect 29929 16949 29963 16983
rect 6009 16745 6043 16779
rect 9413 16677 9447 16711
rect 9781 16677 9815 16711
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 8493 16609 8527 16643
rect 10701 16609 10735 16643
rect 11713 16609 11747 16643
rect 11897 16609 11931 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 15485 16609 15519 16643
rect 15669 16609 15703 16643
rect 16773 16609 16807 16643
rect 19717 16609 19751 16643
rect 22477 16609 22511 16643
rect 22661 16609 22695 16643
rect 23765 16609 23799 16643
rect 25237 16609 25271 16643
rect 25789 16609 25823 16643
rect 27077 16609 27111 16643
rect 27261 16609 27295 16643
rect 28457 16609 28491 16643
rect 1777 16541 1811 16575
rect 3985 16541 4019 16575
rect 5917 16541 5951 16575
rect 8309 16541 8343 16575
rect 10425 16541 10459 16575
rect 14565 16541 14599 16575
rect 15393 16541 15427 16575
rect 17601 16541 17635 16575
rect 18245 16541 18279 16575
rect 18705 16541 18739 16575
rect 19441 16541 19475 16575
rect 22385 16541 22419 16575
rect 23673 16541 23707 16575
rect 28181 16541 28215 16575
rect 28273 16541 28307 16575
rect 2513 16473 2547 16507
rect 5181 16473 5215 16507
rect 9229 16473 9263 16507
rect 13369 16473 13403 16507
rect 21465 16473 21499 16507
rect 26985 16473 27019 16507
rect 6653 16405 6687 16439
rect 7021 16405 7055 16439
rect 7849 16405 7883 16439
rect 8217 16405 8251 16439
rect 10057 16405 10091 16439
rect 10517 16405 10551 16439
rect 11253 16405 11287 16439
rect 11621 16405 11655 16439
rect 12265 16405 12299 16439
rect 13001 16405 13035 16439
rect 14381 16405 14415 16439
rect 15025 16405 15059 16439
rect 17417 16405 17451 16439
rect 18061 16405 18095 16439
rect 22017 16405 22051 16439
rect 23213 16405 23247 16439
rect 23581 16405 23615 16439
rect 24685 16405 24719 16439
rect 25053 16405 25087 16439
rect 25145 16405 25179 16439
rect 25881 16405 25915 16439
rect 26617 16405 26651 16439
rect 27813 16405 27847 16439
rect 7297 16201 7331 16235
rect 10241 16201 10275 16235
rect 23765 16201 23799 16235
rect 24501 16201 24535 16235
rect 26617 16201 26651 16235
rect 26985 16201 27019 16235
rect 27721 16201 27755 16235
rect 4353 16133 4387 16167
rect 8769 16133 8803 16167
rect 10609 16133 10643 16167
rect 12265 16133 12299 16167
rect 19717 16133 19751 16167
rect 20453 16133 20487 16167
rect 23673 16133 23707 16167
rect 24409 16133 24443 16167
rect 1777 16065 1811 16099
rect 3525 16065 3559 16099
rect 5641 16065 5675 16099
rect 7665 16065 7699 16099
rect 8493 16065 8527 16099
rect 11161 16065 11195 16099
rect 11989 16065 12023 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 16313 16065 16347 16099
rect 17785 16065 17819 16099
rect 17877 16065 17911 16099
rect 18613 16065 18647 16099
rect 20545 16065 20579 16099
rect 21465 16049 21499 16083
rect 22293 16065 22327 16099
rect 24869 16065 24903 16099
rect 2053 15997 2087 16031
rect 5733 15997 5767 16031
rect 5917 15997 5951 16031
rect 6653 15997 6687 16031
rect 7757 15997 7791 16031
rect 7941 15997 7975 16031
rect 14841 15997 14875 16031
rect 15485 15997 15519 16031
rect 17969 15997 18003 16031
rect 18889 15997 18923 16031
rect 20729 15997 20763 16031
rect 22017 15997 22051 16031
rect 23949 15997 23983 16031
rect 25145 15997 25179 16031
rect 5273 15929 5307 15963
rect 10977 15929 11011 15963
rect 16681 15929 16715 15963
rect 17417 15929 17451 15963
rect 20085 15929 20119 15963
rect 13737 15861 13771 15895
rect 14289 15861 14323 15895
rect 16129 15861 16163 15895
rect 16957 15861 16991 15895
rect 21281 15861 21315 15895
rect 23305 15861 23339 15895
rect 7849 15657 7883 15691
rect 9321 15657 9355 15691
rect 13185 15657 13219 15691
rect 24501 15657 24535 15691
rect 12081 15589 12115 15623
rect 13553 15589 13587 15623
rect 14473 15589 14507 15623
rect 15853 15589 15887 15623
rect 22753 15589 22787 15623
rect 2053 15521 2087 15555
rect 4629 15521 4663 15555
rect 5641 15521 5675 15555
rect 5825 15521 5859 15555
rect 6837 15521 6871 15555
rect 6929 15521 6963 15555
rect 8401 15521 8435 15555
rect 11437 15521 11471 15555
rect 12725 15521 12759 15555
rect 15025 15521 15059 15555
rect 16497 15521 16531 15555
rect 17049 15521 17083 15555
rect 20269 15521 20303 15555
rect 25789 15521 25823 15555
rect 1777 15453 1811 15487
rect 12449 15453 12483 15487
rect 13737 15453 13771 15487
rect 14841 15453 14875 15487
rect 19625 15453 19659 15487
rect 22293 15453 22327 15487
rect 23121 15453 23155 15487
rect 5549 15385 5583 15419
rect 6745 15385 6779 15419
rect 8309 15385 8343 15419
rect 9229 15385 9263 15419
rect 9781 15385 9815 15419
rect 9965 15385 9999 15419
rect 10241 15385 10275 15419
rect 11253 15385 11287 15419
rect 15485 15385 15519 15419
rect 16221 15385 16255 15419
rect 17325 15385 17359 15419
rect 20545 15385 20579 15419
rect 23949 15385 23983 15419
rect 26249 15385 26283 15419
rect 3985 15317 4019 15351
rect 4353 15317 4387 15351
rect 4445 15317 4479 15351
rect 5181 15317 5215 15351
rect 6377 15317 6411 15351
rect 7481 15317 7515 15351
rect 8217 15317 8251 15351
rect 10885 15317 10919 15351
rect 11345 15317 11379 15351
rect 12541 15317 12575 15351
rect 14197 15317 14231 15351
rect 14933 15317 14967 15351
rect 16313 15317 16347 15351
rect 18797 15317 18831 15351
rect 19441 15317 19475 15351
rect 22017 15317 22051 15351
rect 25237 15317 25271 15351
rect 25605 15317 25639 15351
rect 25697 15317 25731 15351
rect 26433 15317 26467 15351
rect 3525 15113 3559 15147
rect 6745 15113 6779 15147
rect 9597 15113 9631 15147
rect 13001 15113 13035 15147
rect 18429 15113 18463 15147
rect 23765 15113 23799 15147
rect 24041 15113 24075 15147
rect 24225 15113 24259 15147
rect 26985 15113 27019 15147
rect 4445 15045 4479 15079
rect 7665 15045 7699 15079
rect 8585 15045 8619 15079
rect 8769 15045 8803 15079
rect 9689 15045 9723 15079
rect 10793 15045 10827 15079
rect 13461 15045 13495 15079
rect 14105 15045 14139 15079
rect 14841 15045 14875 15079
rect 16773 15045 16807 15079
rect 20177 15045 20211 15079
rect 25145 15045 25179 15079
rect 1777 14977 1811 15011
rect 3709 14977 3743 15011
rect 4169 14977 4203 15011
rect 6653 14977 6687 15011
rect 10885 14977 10919 15011
rect 11713 14977 11747 15011
rect 11989 14977 12023 15011
rect 13369 14977 13403 15011
rect 17141 14977 17175 15011
rect 20085 14977 20119 15011
rect 22017 14977 22051 15011
rect 24869 14977 24903 15011
rect 2053 14909 2087 14943
rect 7757 14909 7791 14943
rect 7849 14909 7883 14943
rect 9873 14909 9907 14943
rect 10977 14909 11011 14943
rect 13553 14909 13587 14943
rect 14565 14909 14599 14943
rect 20361 14909 20395 14943
rect 20913 14909 20947 14943
rect 22293 14909 22327 14943
rect 9229 14841 9263 14875
rect 19717 14841 19751 14875
rect 5917 14773 5951 14807
rect 7297 14773 7331 14807
rect 10425 14773 10459 14807
rect 16313 14773 16347 14807
rect 19165 14773 19199 14807
rect 19349 14773 19383 14807
rect 26617 14773 26651 14807
rect 4261 14569 4295 14603
rect 9413 14569 9447 14603
rect 11621 14569 11655 14603
rect 13737 14569 13771 14603
rect 14381 14569 14415 14603
rect 18613 14569 18647 14603
rect 18889 14569 18923 14603
rect 21741 14569 21775 14603
rect 7205 14501 7239 14535
rect 19441 14501 19475 14535
rect 2053 14433 2087 14467
rect 4813 14433 4847 14467
rect 8493 14433 8527 14467
rect 9965 14433 9999 14467
rect 11161 14433 11195 14467
rect 14105 14433 14139 14467
rect 14933 14433 14967 14467
rect 16865 14433 16899 14467
rect 21097 14433 21131 14467
rect 22293 14433 22327 14467
rect 25145 14433 25179 14467
rect 26341 14433 26375 14467
rect 1777 14365 1811 14399
rect 4629 14365 4663 14399
rect 5457 14365 5491 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 9873 14365 9907 14399
rect 10977 14365 11011 14399
rect 11989 14365 12023 14399
rect 14657 14365 14691 14399
rect 19625 14365 19659 14399
rect 26157 14365 26191 14399
rect 26985 14365 27019 14399
rect 5733 14297 5767 14331
rect 12265 14297 12299 14331
rect 17141 14297 17175 14331
rect 21005 14297 21039 14331
rect 22569 14297 22603 14331
rect 24961 14297 24995 14331
rect 25053 14297 25087 14331
rect 4721 14229 4755 14263
rect 7849 14229 7883 14263
rect 8953 14229 8987 14263
rect 9781 14229 9815 14263
rect 10609 14229 10643 14263
rect 11069 14229 11103 14263
rect 16405 14229 16439 14263
rect 20545 14229 20579 14263
rect 20913 14229 20947 14263
rect 21649 14229 21683 14263
rect 24041 14229 24075 14263
rect 24593 14229 24627 14263
rect 25789 14229 25823 14263
rect 26249 14229 26283 14263
rect 26801 14229 26835 14263
rect 3433 14025 3467 14059
rect 4077 14025 4111 14059
rect 4445 14025 4479 14059
rect 5641 14025 5675 14059
rect 6929 14025 6963 14059
rect 7297 14025 7331 14059
rect 7389 14025 7423 14059
rect 8125 14025 8159 14059
rect 11621 14025 11655 14059
rect 11989 14025 12023 14059
rect 12357 14025 12391 14059
rect 13185 14025 13219 14059
rect 14749 14025 14783 14059
rect 15577 14025 15611 14059
rect 18889 14025 18923 14059
rect 19441 14025 19475 14059
rect 20085 14025 20119 14059
rect 23397 14025 23431 14059
rect 24961 14025 24995 14059
rect 5733 13957 5767 13991
rect 8493 13957 8527 13991
rect 8585 13957 8619 13991
rect 13645 13957 13679 13991
rect 15945 13957 15979 13991
rect 21925 13957 21959 13991
rect 25053 13957 25087 13991
rect 25605 13957 25639 13991
rect 25881 13957 25915 13991
rect 1777 13889 1811 13923
rect 3617 13889 3651 13923
rect 6377 13889 6411 13923
rect 6561 13889 6595 13923
rect 13553 13889 13587 13923
rect 16037 13889 16071 13923
rect 17141 13889 17175 13923
rect 19625 13889 19659 13923
rect 20453 13889 20487 13923
rect 20545 13889 20579 13923
rect 22569 13889 22603 13923
rect 22661 13889 22695 13923
rect 23765 13889 23799 13923
rect 25973 13889 26007 13923
rect 2053 13821 2087 13855
rect 4537 13821 4571 13855
rect 4721 13821 4755 13855
rect 5825 13821 5859 13855
rect 7573 13821 7607 13855
rect 8677 13821 8711 13855
rect 9321 13821 9355 13855
rect 11069 13821 11103 13855
rect 12449 13821 12483 13855
rect 12541 13821 12575 13855
rect 13829 13821 13863 13855
rect 14841 13821 14875 13855
rect 15025 13821 15059 13855
rect 16221 13821 16255 13855
rect 17417 13821 17451 13855
rect 20637 13821 20671 13855
rect 22845 13821 22879 13855
rect 23857 13821 23891 13855
rect 24041 13821 24075 13855
rect 25145 13821 25179 13855
rect 14381 13753 14415 13787
rect 22201 13753 22235 13787
rect 5273 13685 5307 13719
rect 9584 13685 9618 13719
rect 16681 13685 16715 13719
rect 24593 13685 24627 13719
rect 6285 13481 6319 13515
rect 11621 13481 11655 13515
rect 13737 13481 13771 13515
rect 16037 13481 16071 13515
rect 18889 13481 18923 13515
rect 22109 13481 22143 13515
rect 23949 13481 23983 13515
rect 11437 13413 11471 13447
rect 22845 13413 22879 13447
rect 24133 13413 24167 13447
rect 2789 13345 2823 13379
rect 4169 13345 4203 13379
rect 6745 13345 6779 13379
rect 9137 13345 9171 13379
rect 9413 13345 9447 13379
rect 10977 13345 11011 13379
rect 11989 13345 12023 13379
rect 14565 13345 14599 13379
rect 17141 13345 17175 13379
rect 20361 13345 20395 13379
rect 23305 13345 23339 13379
rect 23489 13345 23523 13379
rect 1777 13277 1811 13311
rect 14289 13277 14323 13311
rect 22477 13277 22511 13311
rect 3341 13209 3375 13243
rect 4445 13209 4479 13243
rect 7021 13209 7055 13243
rect 10885 13209 10919 13243
rect 12265 13209 12299 13243
rect 17417 13209 17451 13243
rect 20637 13209 20671 13243
rect 23213 13209 23247 13243
rect 24593 13209 24627 13243
rect 25421 13209 25455 13243
rect 5917 13141 5951 13175
rect 8493 13141 8527 13175
rect 10425 13141 10459 13175
rect 10793 13141 10827 13175
rect 16497 13141 16531 13175
rect 19349 13141 19383 13175
rect 19441 13141 19475 13175
rect 4997 12937 5031 12971
rect 5733 12937 5767 12971
rect 7297 12937 7331 12971
rect 10517 12937 10551 12971
rect 10977 12937 11011 12971
rect 12541 12937 12575 12971
rect 17785 12937 17819 12971
rect 18153 12937 18187 12971
rect 21097 12937 21131 12971
rect 22201 12937 22235 12971
rect 24777 12937 24811 12971
rect 3709 12869 3743 12903
rect 4261 12869 4295 12903
rect 5641 12869 5675 12903
rect 11897 12869 11931 12903
rect 14105 12869 14139 12903
rect 15669 12869 15703 12903
rect 16405 12869 16439 12903
rect 18981 12869 19015 12903
rect 1593 12801 1627 12835
rect 2697 12801 2731 12835
rect 3525 12801 3559 12835
rect 7205 12801 7239 12835
rect 10057 12801 10091 12835
rect 10701 12801 10735 12835
rect 12909 12801 12943 12835
rect 14933 12801 14967 12835
rect 18245 12801 18279 12835
rect 21189 12801 21223 12835
rect 23029 12801 23063 12835
rect 1869 12733 1903 12767
rect 5917 12733 5951 12767
rect 7389 12733 7423 12767
rect 8033 12733 8067 12767
rect 8309 12733 8343 12767
rect 13001 12733 13035 12767
rect 13093 12733 13127 12767
rect 14197 12733 14231 12767
rect 14381 12733 14415 12767
rect 16865 12733 16899 12767
rect 18429 12733 18463 12767
rect 19809 12733 19843 12767
rect 21373 12733 21407 12767
rect 23305 12733 23339 12767
rect 4445 12665 4479 12699
rect 11253 12665 11287 12699
rect 5273 12597 5307 12631
rect 6837 12597 6871 12631
rect 11621 12597 11655 12631
rect 13737 12597 13771 12631
rect 16129 12597 16163 12631
rect 20729 12597 20763 12631
rect 25053 12597 25087 12631
rect 3065 12393 3099 12427
rect 3985 12393 4019 12427
rect 4629 12393 4663 12427
rect 7849 12393 7883 12427
rect 11805 12393 11839 12427
rect 14197 12393 14231 12427
rect 14381 12393 14415 12427
rect 18061 12393 18095 12427
rect 21833 12393 21867 12427
rect 24409 12393 24443 12427
rect 1869 12257 1903 12291
rect 4721 12257 4755 12291
rect 5365 12257 5399 12291
rect 7389 12257 7423 12291
rect 8401 12257 8435 12291
rect 9873 12257 9907 12291
rect 11253 12257 11287 12291
rect 12357 12257 12391 12291
rect 13645 12257 13679 12291
rect 16589 12257 16623 12291
rect 18337 12257 18371 12291
rect 20085 12257 20119 12291
rect 20361 12257 20395 12291
rect 22569 12257 22603 12291
rect 1593 12189 1627 12223
rect 2973 12189 3007 12223
rect 3433 12189 3467 12223
rect 3893 12189 3927 12223
rect 4169 12189 4203 12223
rect 8309 12189 8343 12223
rect 11069 12189 11103 12223
rect 12173 12189 12207 12223
rect 13369 12189 13403 12223
rect 14749 12189 14783 12223
rect 15945 12189 15979 12223
rect 16313 12189 16347 12223
rect 19533 12189 19567 12223
rect 22293 12189 22327 12223
rect 5641 12121 5675 12155
rect 9137 12121 9171 12155
rect 15485 12121 15519 12155
rect 18889 12121 18923 12155
rect 8217 12053 8251 12087
rect 10609 12053 10643 12087
rect 10977 12053 11011 12087
rect 12265 12053 12299 12087
rect 13001 12053 13035 12087
rect 13461 12053 13495 12087
rect 18521 12053 18555 12087
rect 18981 12053 19015 12087
rect 19349 12053 19383 12087
rect 24041 12053 24075 12087
rect 1409 11849 1443 11883
rect 4445 11849 4479 11883
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 6745 11849 6779 11883
rect 11713 11849 11747 11883
rect 15209 11849 15243 11883
rect 15577 11849 15611 11883
rect 16037 11849 16071 11883
rect 17417 11849 17451 11883
rect 18153 11849 18187 11883
rect 18613 11849 18647 11883
rect 19349 11849 19383 11883
rect 21925 11849 21959 11883
rect 24409 11849 24443 11883
rect 3341 11781 3375 11815
rect 3433 11781 3467 11815
rect 5733 11781 5767 11815
rect 7665 11781 7699 11815
rect 12449 11781 12483 11815
rect 18521 11781 18555 11815
rect 19165 11781 19199 11815
rect 22661 11781 22695 11815
rect 2421 11713 2455 11747
rect 4537 11713 4571 11747
rect 7389 11713 7423 11747
rect 9597 11713 9631 11747
rect 12357 11713 12391 11747
rect 13185 11713 13219 11747
rect 15945 11713 15979 11747
rect 17325 11713 17359 11747
rect 2145 11645 2179 11679
rect 4721 11645 4755 11679
rect 5917 11645 5951 11679
rect 10333 11645 10367 11679
rect 10977 11645 11011 11679
rect 12541 11645 12575 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 17601 11645 17635 11679
rect 18705 11645 18739 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 22385 11645 22419 11679
rect 9137 11577 9171 11611
rect 4077 11509 4111 11543
rect 11989 11509 12023 11543
rect 14933 11509 14967 11543
rect 16957 11509 16991 11543
rect 21465 11509 21499 11543
rect 24133 11509 24167 11543
rect 5076 11305 5110 11339
rect 6561 11305 6595 11339
rect 13645 11305 13679 11339
rect 16497 11305 16531 11339
rect 18889 11305 18923 11339
rect 22661 11305 22695 11339
rect 23029 11305 23063 11339
rect 32045 11305 32079 11339
rect 4261 11237 4295 11271
rect 7849 11237 7883 11271
rect 2237 11169 2271 11203
rect 2513 11169 2547 11203
rect 3617 11169 3651 11203
rect 4813 11169 4847 11203
rect 8401 11169 8435 11203
rect 9597 11169 9631 11203
rect 9689 11169 9723 11203
rect 10977 11169 11011 11203
rect 11529 11169 11563 11203
rect 13277 11169 13311 11203
rect 29745 11169 29779 11203
rect 1777 11101 1811 11135
rect 3433 11101 3467 11135
rect 7021 11101 7055 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 14749 11101 14783 11135
rect 17141 11101 17175 11135
rect 19533 11101 19567 11135
rect 20913 11101 20947 11135
rect 31769 11101 31803 11135
rect 4077 11033 4111 11067
rect 10701 11033 10735 11067
rect 11805 11033 11839 11067
rect 15025 11033 15059 11067
rect 17417 11033 17451 11067
rect 20269 11033 20303 11067
rect 21189 11033 21223 11067
rect 30021 11033 30055 11067
rect 1593 10965 1627 10999
rect 7481 10965 7515 10999
rect 8309 10965 8343 10999
rect 9137 10965 9171 10999
rect 10333 10965 10367 10999
rect 10793 10965 10827 10999
rect 16773 10965 16807 10999
rect 5825 10761 5859 10795
rect 9965 10761 9999 10795
rect 10793 10761 10827 10795
rect 13829 10761 13863 10795
rect 14381 10761 14415 10795
rect 14841 10761 14875 10795
rect 19257 10761 19291 10795
rect 21833 10761 21867 10795
rect 22017 10761 22051 10795
rect 6561 10693 6595 10727
rect 10701 10693 10735 10727
rect 12357 10693 12391 10727
rect 17785 10693 17819 10727
rect 2145 10625 2179 10659
rect 2421 10625 2455 10659
rect 3433 10625 3467 10659
rect 5365 10625 5399 10659
rect 7021 10625 7055 10659
rect 14749 10625 14783 10659
rect 15945 10625 15979 10659
rect 17509 10625 17543 10659
rect 3709 10557 3743 10591
rect 7481 10557 7515 10591
rect 7757 10557 7791 10591
rect 9505 10557 9539 10591
rect 10885 10557 10919 10591
rect 12081 10557 12115 10591
rect 15025 10557 15059 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 16865 10557 16899 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 10333 10489 10367 10523
rect 15577 10489 15611 10523
rect 5181 10421 5215 10455
rect 6837 10421 6871 10455
rect 9781 10421 9815 10455
rect 11529 10421 11563 10455
rect 21465 10421 21499 10455
rect 3249 10217 3283 10251
rect 6561 10217 6595 10251
rect 9045 10217 9079 10251
rect 10057 10217 10091 10251
rect 8585 10149 8619 10183
rect 14105 10149 14139 10183
rect 18889 10149 18923 10183
rect 21557 10149 21591 10183
rect 1593 10081 1627 10115
rect 1869 10081 1903 10115
rect 4537 10081 4571 10115
rect 5825 10081 5859 10115
rect 6837 10081 6871 10115
rect 10517 10081 10551 10115
rect 10701 10081 10735 10115
rect 13553 10081 13587 10115
rect 14841 10081 14875 10115
rect 19441 10081 19475 10115
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 4261 10013 4295 10047
rect 9413 10013 9447 10047
rect 11253 10013 11287 10047
rect 14565 10013 14599 10047
rect 17141 10013 17175 10047
rect 3985 9945 4019 9979
rect 7113 9945 7147 9979
rect 11529 9945 11563 9979
rect 17417 9945 17451 9979
rect 19717 9945 19751 9979
rect 10425 9877 10459 9911
rect 13001 9877 13035 9911
rect 16313 9877 16347 9911
rect 16589 9877 16623 9911
rect 16773 9877 16807 9911
rect 21189 9877 21223 9911
rect 1501 9673 1535 9707
rect 13829 9673 13863 9707
rect 13921 9673 13955 9707
rect 16221 9673 16255 9707
rect 1593 9605 1627 9639
rect 5733 9605 5767 9639
rect 5825 9605 5859 9639
rect 8401 9605 8435 9639
rect 11989 9605 12023 9639
rect 17141 9605 17175 9639
rect 19533 9605 19567 9639
rect 28457 9605 28491 9639
rect 2237 9537 2271 9571
rect 3801 9537 3835 9571
rect 4261 9537 4295 9571
rect 7113 9537 7147 9571
rect 8132 9537 8166 9571
rect 10701 9537 10735 9571
rect 19441 9537 19475 9571
rect 27537 9537 27571 9571
rect 1961 9469 1995 9503
rect 4537 9469 4571 9503
rect 6745 9469 6779 9503
rect 6837 9469 6871 9503
rect 10793 9469 10827 9503
rect 10885 9469 10919 9503
rect 11713 9469 11747 9503
rect 14473 9469 14507 9503
rect 14749 9469 14783 9503
rect 16865 9469 16899 9503
rect 19717 9469 19751 9503
rect 27997 9469 28031 9503
rect 3617 9401 3651 9435
rect 19073 9401 19107 9435
rect 9873 9333 9907 9367
rect 10333 9333 10367 9367
rect 13461 9333 13495 9367
rect 18613 9333 18647 9367
rect 20085 9333 20119 9367
rect 27813 9333 27847 9367
rect 3801 9129 3835 9163
rect 4629 9129 4663 9163
rect 7205 9129 7239 9163
rect 7849 9129 7883 9163
rect 10149 9129 10183 9163
rect 11575 9129 11609 9163
rect 14289 9061 14323 9095
rect 1593 8993 1627 9027
rect 1869 8993 1903 9027
rect 3985 8993 4019 9027
rect 4721 8993 4755 9027
rect 6193 8993 6227 9027
rect 8401 8993 8435 9027
rect 9413 8993 9447 9027
rect 10793 8993 10827 9027
rect 14933 8993 14967 9027
rect 16037 8993 16071 9027
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 5917 8925 5951 8959
rect 7389 8925 7423 8959
rect 8217 8925 8251 8959
rect 11345 8925 11379 8959
rect 14749 8925 14783 8959
rect 10517 8857 10551 8891
rect 13553 8857 13587 8891
rect 14657 8857 14691 8891
rect 16313 8857 16347 8891
rect 2881 8789 2915 8823
rect 8309 8789 8343 8823
rect 9045 8789 9079 8823
rect 10609 8789 10643 8823
rect 12633 8789 12667 8823
rect 17785 8789 17819 8823
rect 18153 8789 18187 8823
rect 18705 8789 18739 8823
rect 18981 8789 19015 8823
rect 3341 8585 3375 8619
rect 3985 8585 4019 8619
rect 5825 8585 5859 8619
rect 7297 8585 7331 8619
rect 10149 8585 10183 8619
rect 12541 8585 12575 8619
rect 14289 8585 14323 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 3525 8517 3559 8551
rect 5181 8517 5215 8551
rect 7205 8517 7239 8551
rect 1593 8449 1627 8483
rect 3065 8449 3099 8483
rect 4169 8449 4203 8483
rect 4813 8449 4847 8483
rect 6009 8449 6043 8483
rect 7757 8449 7791 8483
rect 8677 8449 8711 8483
rect 10517 8449 10551 8483
rect 13645 8449 13679 8483
rect 14657 8449 14691 8483
rect 1869 8381 1903 8415
rect 8401 8381 8435 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 12633 8381 12667 8415
rect 12817 8381 12851 8415
rect 14749 8381 14783 8415
rect 14933 8381 14967 8415
rect 16037 8381 16071 8415
rect 16221 8381 16255 8415
rect 2881 8313 2915 8347
rect 4629 8313 4663 8347
rect 9597 8313 9631 8347
rect 12173 8313 12207 8347
rect 1593 8041 1627 8075
rect 3801 8041 3835 8075
rect 4353 8041 4387 8075
rect 9597 8041 9631 8075
rect 13001 8041 13035 8075
rect 2881 7973 2915 8007
rect 15209 7973 15243 8007
rect 3525 7905 3559 7939
rect 10057 7905 10091 7939
rect 10149 7905 10183 7939
rect 11529 7905 11563 7939
rect 13553 7905 13587 7939
rect 14841 7905 14875 7939
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 3341 7837 3375 7871
rect 11253 7837 11287 7871
rect 13461 7837 13495 7871
rect 15025 7837 15059 7871
rect 11161 7769 11195 7803
rect 2237 7701 2271 7735
rect 9965 7701 9999 7735
rect 13369 7701 13403 7735
rect 1593 7497 1627 7531
rect 2237 7497 2271 7531
rect 3525 7497 3559 7531
rect 9137 7497 9171 7531
rect 11897 7497 11931 7531
rect 13461 7497 13495 7531
rect 23949 7497 23983 7531
rect 4169 7429 4203 7463
rect 24225 7429 24259 7463
rect 1777 7361 1811 7395
rect 2421 7361 2455 7395
rect 3065 7361 3099 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 9321 7361 9355 7395
rect 10793 7361 10827 7395
rect 12725 7361 12759 7395
rect 14289 7361 14323 7395
rect 22201 7361 22235 7395
rect 4353 7293 4387 7327
rect 22477 7293 22511 7327
rect 10609 7225 10643 7259
rect 2881 7157 2915 7191
rect 12541 7157 12575 7191
rect 14105 7157 14139 7191
rect 2237 6953 2271 6987
rect 23213 6953 23247 6987
rect 3341 6885 3375 6919
rect 3801 6817 3835 6851
rect 10609 6817 10643 6851
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 3525 6749 3559 6783
rect 22937 6749 22971 6783
rect 1593 6613 1627 6647
rect 2881 6613 2915 6647
rect 3985 6613 4019 6647
rect 23397 6613 23431 6647
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 22452 6273 22486 6307
rect 1593 6205 1627 6239
rect 1869 6205 1903 6239
rect 2881 6137 2915 6171
rect 22523 6069 22557 6103
rect 2697 5865 2731 5899
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 15577 5729 15611 5763
rect 15761 5729 15795 5763
rect 17141 5729 17175 5763
rect 24869 5729 24903 5763
rect 26985 5729 27019 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 20913 5661 20947 5695
rect 24685 5661 24719 5695
rect 2881 5593 2915 5627
rect 17417 5593 17451 5627
rect 19349 5593 19383 5627
rect 26525 5593 26559 5627
rect 27169 5593 27203 5627
rect 28825 5593 28859 5627
rect 16221 5525 16255 5559
rect 21373 5525 21407 5559
rect 22891 5321 22925 5355
rect 1593 5185 1627 5219
rect 2697 5185 2731 5219
rect 15669 5185 15703 5219
rect 17509 5185 17543 5219
rect 22144 5185 22178 5219
rect 22788 5185 22822 5219
rect 1869 5117 1903 5151
rect 15853 5117 15887 5151
rect 17693 5117 17727 5151
rect 28641 5117 28675 5151
rect 28825 5117 28859 5151
rect 30297 5117 30331 5151
rect 16313 4981 16347 5015
rect 18153 4981 18187 5015
rect 22247 4981 22281 5015
rect 19533 4777 19567 4811
rect 24731 4777 24765 4811
rect 1593 4641 1627 4675
rect 1869 4641 1903 4675
rect 25973 4641 26007 4675
rect 27537 4641 27571 4675
rect 2881 4573 2915 4607
rect 19441 4573 19475 4607
rect 24628 4573 24662 4607
rect 25789 4573 25823 4607
rect 2789 4437 2823 4471
rect 19901 4437 19935 4471
rect 2237 4233 2271 4267
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 3065 4097 3099 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 15209 4097 15243 4131
rect 2881 3961 2915 3995
rect 1593 3893 1627 3927
rect 15025 3893 15059 3927
rect 2881 3689 2915 3723
rect 3525 3621 3559 3655
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 11529 3485 11563 3519
rect 1823 3349 1857 3383
rect 3341 3349 3375 3383
rect 11621 3349 11655 3383
rect 2881 3145 2915 3179
rect 12725 3145 12759 3179
rect 12633 3077 12667 3111
rect 13921 3077 13955 3111
rect 15577 3077 15611 3111
rect 1869 3009 1903 3043
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 8769 3009 8803 3043
rect 17049 3009 17083 3043
rect 18337 3009 18371 3043
rect 20545 3009 20579 3043
rect 1593 2941 1627 2975
rect 3525 2941 3559 2975
rect 9045 2941 9079 2975
rect 14105 2941 14139 2975
rect 10517 2873 10551 2907
rect 15761 2873 15795 2907
rect 10793 2805 10827 2839
rect 16865 2805 16899 2839
rect 18153 2805 18187 2839
rect 20361 2805 20395 2839
rect 2881 2601 2915 2635
rect 25513 2601 25547 2635
rect 28181 2601 28215 2635
rect 30849 2601 30883 2635
rect 33517 2601 33551 2635
rect 1593 2465 1627 2499
rect 3525 2465 3559 2499
rect 4629 2465 4663 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 15301 2465 15335 2499
rect 17969 2465 18003 2499
rect 20545 2465 20579 2499
rect 23121 2465 23155 2499
rect 36369 2465 36403 2499
rect 1869 2397 1903 2431
rect 3065 2397 3099 2431
rect 3341 2397 3375 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17509 2397 17543 2431
rect 20085 2397 20119 2431
rect 22661 2397 22695 2431
rect 25697 2397 25731 2431
rect 25973 2397 26007 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33701 2397 33735 2431
rect 33977 2397 34011 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
<< metal1 >>
rect 22830 25644 22836 25696
rect 22888 25684 22894 25696
rect 27798 25684 27804 25696
rect 22888 25656 27804 25684
rect 22888 25644 22894 25656
rect 27798 25644 27804 25656
rect 27856 25644 27862 25696
rect 10134 25576 10140 25628
rect 10192 25616 10198 25628
rect 33594 25616 33600 25628
rect 10192 25588 33600 25616
rect 10192 25576 10198 25588
rect 33594 25576 33600 25588
rect 33652 25576 33658 25628
rect 7006 25508 7012 25560
rect 7064 25548 7070 25560
rect 32858 25548 32864 25560
rect 7064 25520 32864 25548
rect 7064 25508 7070 25520
rect 32858 25508 32864 25520
rect 32916 25508 32922 25560
rect 10870 25440 10876 25492
rect 10928 25480 10934 25492
rect 35618 25480 35624 25492
rect 10928 25452 35624 25480
rect 10928 25440 10934 25452
rect 35618 25440 35624 25452
rect 35676 25440 35682 25492
rect 15838 25372 15844 25424
rect 15896 25412 15902 25424
rect 34238 25412 34244 25424
rect 15896 25384 34244 25412
rect 15896 25372 15902 25384
rect 34238 25372 34244 25384
rect 34296 25372 34302 25424
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 31570 25344 31576 25356
rect 10100 25316 31576 25344
rect 10100 25304 10106 25316
rect 31570 25304 31576 25316
rect 31628 25304 31634 25356
rect 12066 25236 12072 25288
rect 12124 25276 12130 25288
rect 33778 25276 33784 25288
rect 12124 25248 33784 25276
rect 12124 25236 12130 25248
rect 33778 25236 33784 25248
rect 33836 25236 33842 25288
rect 12618 25168 12624 25220
rect 12676 25208 12682 25220
rect 34790 25208 34796 25220
rect 12676 25180 34796 25208
rect 12676 25168 12682 25180
rect 34790 25168 34796 25180
rect 34848 25168 34854 25220
rect 9858 25100 9864 25152
rect 9916 25140 9922 25152
rect 31754 25140 31760 25152
rect 9916 25112 31760 25140
rect 9916 25100 9922 25112
rect 31754 25100 31760 25112
rect 31812 25100 31818 25152
rect 10778 25032 10784 25084
rect 10836 25072 10842 25084
rect 34606 25072 34612 25084
rect 10836 25044 34612 25072
rect 10836 25032 10842 25044
rect 34606 25032 34612 25044
rect 34664 25032 34670 25084
rect 14918 24964 14924 25016
rect 14976 25004 14982 25016
rect 31110 25004 31116 25016
rect 14976 24976 31116 25004
rect 14976 24964 14982 24976
rect 31110 24964 31116 24976
rect 31168 24964 31174 25016
rect 4062 24896 4068 24948
rect 4120 24936 4126 24948
rect 7466 24936 7472 24948
rect 4120 24908 7472 24936
rect 4120 24896 4126 24908
rect 7466 24896 7472 24908
rect 7524 24896 7530 24948
rect 15378 24896 15384 24948
rect 15436 24936 15442 24948
rect 33686 24936 33692 24948
rect 15436 24908 33692 24936
rect 15436 24896 15442 24908
rect 33686 24896 33692 24908
rect 33744 24896 33750 24948
rect 12802 24828 12808 24880
rect 12860 24868 12866 24880
rect 32030 24868 32036 24880
rect 12860 24840 32036 24868
rect 12860 24828 12866 24840
rect 32030 24828 32036 24840
rect 32088 24828 32094 24880
rect 11698 24760 11704 24812
rect 11756 24800 11762 24812
rect 22002 24800 22008 24812
rect 11756 24772 22008 24800
rect 11756 24760 11762 24772
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 22554 24760 22560 24812
rect 22612 24800 22618 24812
rect 30006 24800 30012 24812
rect 22612 24772 30012 24800
rect 22612 24760 22618 24772
rect 30006 24760 30012 24772
rect 30064 24760 30070 24812
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 26050 24732 26056 24744
rect 14332 24704 26056 24732
rect 14332 24692 14338 24704
rect 26050 24692 26056 24704
rect 26108 24692 26114 24744
rect 30374 24732 30380 24744
rect 28184 24704 30380 24732
rect 12342 24624 12348 24676
rect 12400 24664 12406 24676
rect 25774 24664 25780 24676
rect 12400 24636 25780 24664
rect 12400 24624 12406 24636
rect 25774 24624 25780 24636
rect 25832 24624 25838 24676
rect 25958 24624 25964 24676
rect 26016 24664 26022 24676
rect 28184 24664 28212 24704
rect 30374 24692 30380 24704
rect 30432 24692 30438 24744
rect 26016 24636 28212 24664
rect 26016 24624 26022 24636
rect 28258 24624 28264 24676
rect 28316 24664 28322 24676
rect 31202 24664 31208 24676
rect 28316 24636 31208 24664
rect 28316 24624 28322 24636
rect 31202 24624 31208 24636
rect 31260 24624 31266 24676
rect 35894 24624 35900 24676
rect 35952 24664 35958 24676
rect 36814 24664 36820 24676
rect 35952 24636 36820 24664
rect 35952 24624 35958 24636
rect 36814 24624 36820 24636
rect 36872 24624 36878 24676
rect 17126 24556 17132 24608
rect 17184 24596 17190 24608
rect 18782 24596 18788 24608
rect 17184 24568 18788 24596
rect 17184 24556 17190 24568
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 25130 24556 25136 24608
rect 25188 24596 25194 24608
rect 28994 24596 29000 24608
rect 25188 24568 29000 24596
rect 25188 24556 25194 24568
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 29086 24556 29092 24608
rect 29144 24596 29150 24608
rect 40310 24596 40316 24608
rect 29144 24568 40316 24596
rect 29144 24556 29150 24568
rect 40310 24556 40316 24568
rect 40368 24556 40374 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 3973 24395 4031 24401
rect 3973 24361 3985 24395
rect 4019 24392 4031 24395
rect 4019 24364 11652 24392
rect 4019 24361 4031 24364
rect 3973 24355 4031 24361
rect 2038 24284 2044 24336
rect 2096 24324 2102 24336
rect 9306 24324 9312 24336
rect 2096 24296 4660 24324
rect 2096 24284 2102 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2314 24188 2320 24200
rect 2271 24160 2320 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4246 24188 4252 24200
rect 4203 24160 4252 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4246 24148 4252 24160
rect 4304 24148 4310 24200
rect 4632 24197 4660 24296
rect 8220 24296 9312 24324
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 7098 24256 7104 24268
rect 5859 24228 7104 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 7098 24216 7104 24228
rect 7156 24216 7162 24268
rect 8220 24265 8248 24296
rect 9306 24284 9312 24296
rect 9364 24284 9370 24336
rect 11624 24324 11652 24364
rect 11698 24352 11704 24404
rect 11756 24352 11762 24404
rect 14274 24352 14280 24404
rect 14332 24352 14338 24404
rect 18966 24392 18972 24404
rect 16776 24364 18972 24392
rect 14458 24324 14464 24336
rect 11624 24296 12434 24324
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24225 8263 24259
rect 8205 24219 8263 24225
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 12406 24256 12434 24296
rect 13556 24296 14464 24324
rect 13556 24265 13584 24296
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 13541 24259 13599 24265
rect 11011 24228 12020 24256
rect 12406 24228 13216 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 6638 24148 6644 24200
rect 6696 24188 6702 24200
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6696 24160 6745 24188
rect 6696 24148 6702 24160
rect 6733 24157 6745 24160
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 7190 24148 7196 24200
rect 7248 24148 7254 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10042 24188 10048 24200
rect 9999 24160 10048 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 3602 24012 3608 24064
rect 3660 24052 3666 24064
rect 5994 24052 6000 24064
rect 3660 24024 6000 24052
rect 3660 24012 3666 24024
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 6546 24012 6552 24064
rect 6604 24012 6610 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 9324 24052 9352 24151
rect 10042 24148 10048 24160
rect 10100 24148 10106 24200
rect 11882 24148 11888 24200
rect 11940 24148 11946 24200
rect 11992 24120 12020 24228
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12618 24188 12624 24200
rect 12575 24160 12624 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 13188 24188 13216 24228
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 16776 24256 16804 24364
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 20162 24352 20168 24404
rect 20220 24392 20226 24404
rect 38565 24395 38623 24401
rect 38565 24392 38577 24395
rect 20220 24364 38577 24392
rect 20220 24352 20226 24364
rect 38565 24361 38577 24364
rect 38611 24361 38623 24395
rect 38565 24355 38623 24361
rect 41506 24352 41512 24404
rect 41564 24392 41570 24404
rect 42153 24395 42211 24401
rect 42153 24392 42165 24395
rect 41564 24364 42165 24392
rect 41564 24352 41570 24364
rect 42153 24361 42165 24364
rect 42199 24361 42211 24395
rect 42153 24355 42211 24361
rect 18138 24284 18144 24336
rect 18196 24324 18202 24336
rect 18196 24296 18828 24324
rect 18196 24284 18202 24296
rect 16163 24228 16804 24256
rect 16853 24259 16911 24265
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 18690 24256 18696 24268
rect 16899 24228 18696 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 18800 24256 18828 24296
rect 19058 24284 19064 24336
rect 19116 24324 19122 24336
rect 19116 24296 26464 24324
rect 19116 24284 19122 24296
rect 18800 24228 20208 24256
rect 13906 24188 13912 24200
rect 13188 24160 13912 24188
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24157 15163 24191
rect 15105 24151 15163 24157
rect 13814 24120 13820 24132
rect 11992 24092 13820 24120
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 15120 24120 15148 24151
rect 19518 24148 19524 24200
rect 19576 24188 19582 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 19576 24160 19625 24188
rect 19576 24148 19582 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19886 24148 19892 24200
rect 19944 24188 19950 24200
rect 20073 24191 20131 24197
rect 20073 24188 20085 24191
rect 19944 24160 20085 24188
rect 19944 24148 19950 24160
rect 20073 24157 20085 24160
rect 20119 24157 20131 24191
rect 20180 24188 20208 24228
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 21600 24228 22477 24256
rect 21600 24216 21606 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 25038 24256 25044 24268
rect 22465 24219 22523 24225
rect 24044 24228 25044 24256
rect 21174 24188 21180 24200
rect 20180 24160 21180 24188
rect 20073 24151 20131 24157
rect 21174 24148 21180 24160
rect 21232 24148 21238 24200
rect 22002 24148 22008 24200
rect 22060 24148 22066 24200
rect 22094 24148 22100 24200
rect 22152 24188 22158 24200
rect 24044 24197 24072 24228
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 25130 24216 25136 24268
rect 25188 24216 25194 24268
rect 25222 24216 25228 24268
rect 25280 24256 25286 24268
rect 26329 24259 26387 24265
rect 26329 24256 26341 24259
rect 25280 24228 26341 24256
rect 25280 24216 25286 24228
rect 26329 24225 26341 24228
rect 26375 24225 26387 24259
rect 26436 24256 26464 24296
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 28997 24327 29055 24333
rect 28997 24324 29009 24327
rect 27672 24296 29009 24324
rect 27672 24284 27678 24296
rect 28997 24293 29009 24296
rect 29043 24293 29055 24327
rect 31297 24327 31355 24333
rect 31297 24324 31309 24327
rect 28997 24287 29055 24293
rect 29104 24296 31309 24324
rect 27709 24259 27767 24265
rect 27709 24256 27721 24259
rect 26436 24228 27721 24256
rect 26329 24219 26387 24225
rect 27709 24225 27721 24228
rect 27755 24225 27767 24259
rect 27709 24219 27767 24225
rect 28626 24216 28632 24268
rect 28684 24256 28690 24268
rect 29104 24256 29132 24296
rect 31297 24293 31309 24296
rect 31343 24293 31355 24327
rect 32769 24327 32827 24333
rect 32769 24324 32781 24327
rect 31297 24287 31355 24293
rect 31726 24296 32781 24324
rect 28684 24228 29132 24256
rect 28684 24216 28690 24228
rect 29270 24216 29276 24268
rect 29328 24256 29334 24268
rect 29733 24259 29791 24265
rect 29733 24256 29745 24259
rect 29328 24228 29745 24256
rect 29328 24216 29334 24228
rect 29733 24225 29745 24228
rect 29779 24256 29791 24259
rect 31726 24256 31754 24296
rect 32769 24293 32781 24296
rect 32815 24293 32827 24327
rect 32769 24287 32827 24293
rect 33502 24284 33508 24336
rect 33560 24284 33566 24336
rect 34054 24284 34060 24336
rect 34112 24324 34118 24336
rect 36817 24327 36875 24333
rect 36817 24324 36829 24327
rect 34112 24296 36829 24324
rect 34112 24284 34118 24296
rect 36817 24293 36829 24296
rect 36863 24293 36875 24327
rect 36817 24287 36875 24293
rect 29779 24228 31754 24256
rect 29779 24225 29791 24228
rect 29733 24219 29791 24225
rect 34238 24216 34244 24268
rect 34296 24216 34302 24268
rect 37001 24259 37059 24265
rect 37001 24256 37013 24259
rect 34992 24228 37013 24256
rect 24029 24191 24087 24197
rect 24029 24188 24041 24191
rect 22152 24160 24041 24188
rect 22152 24148 22158 24160
rect 24029 24157 24041 24160
rect 24075 24157 24087 24191
rect 24029 24151 24087 24157
rect 25314 24148 25320 24200
rect 25372 24188 25378 24200
rect 27617 24191 27675 24197
rect 27617 24188 27629 24191
rect 25372 24160 27629 24188
rect 25372 24148 25378 24160
rect 27617 24157 27629 24160
rect 27663 24157 27675 24191
rect 27617 24151 27675 24157
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 17034 24120 17040 24132
rect 15120 24092 17040 24120
rect 17034 24080 17040 24092
rect 17092 24080 17098 24132
rect 17126 24080 17132 24132
rect 17184 24080 17190 24132
rect 18506 24120 18512 24132
rect 18354 24092 18512 24120
rect 18506 24080 18512 24092
rect 18564 24120 18570 24132
rect 18969 24123 19027 24129
rect 18969 24120 18981 24123
rect 18564 24092 18981 24120
rect 18564 24080 18570 24092
rect 18969 24089 18981 24092
rect 19015 24089 19027 24123
rect 25222 24120 25228 24132
rect 18969 24083 19027 24089
rect 19076 24092 25228 24120
rect 13722 24052 13728 24064
rect 9324 24024 13728 24052
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 16942 24012 16948 24064
rect 17000 24052 17006 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 17000 24024 18613 24052
rect 17000 24012 17006 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18601 24015 18659 24021
rect 18782 24012 18788 24064
rect 18840 24052 18846 24064
rect 19076 24052 19104 24092
rect 25222 24080 25228 24092
rect 25280 24080 25286 24132
rect 25958 24120 25964 24132
rect 25700 24092 25964 24120
rect 18840 24024 19104 24052
rect 19429 24055 19487 24061
rect 18840 24012 18846 24024
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 20438 24052 20444 24064
rect 19475 24024 20444 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24052 23903 24055
rect 24486 24052 24492 24064
rect 23891 24024 24492 24052
rect 23891 24021 23903 24024
rect 23845 24015 23903 24021
rect 24486 24012 24492 24024
rect 24544 24012 24550 24064
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 24946 24012 24952 24064
rect 25004 24012 25010 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25700 24052 25728 24092
rect 25958 24080 25964 24092
rect 26016 24080 26022 24132
rect 26050 24080 26056 24132
rect 26108 24120 26114 24132
rect 26237 24123 26295 24129
rect 26237 24120 26249 24123
rect 26108 24092 26249 24120
rect 26108 24080 26114 24092
rect 26237 24089 26249 24092
rect 26283 24089 26295 24123
rect 26237 24083 26295 24089
rect 26694 24080 26700 24132
rect 26752 24120 26758 24132
rect 28552 24120 28580 24151
rect 29178 24148 29184 24200
rect 29236 24148 29242 24200
rect 30006 24148 30012 24200
rect 30064 24148 30070 24200
rect 30558 24148 30564 24200
rect 30616 24188 30622 24200
rect 31478 24188 31484 24200
rect 30616 24160 31484 24188
rect 30616 24148 30622 24160
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 31846 24148 31852 24200
rect 31904 24188 31910 24200
rect 32490 24188 32496 24200
rect 31904 24160 32496 24188
rect 31904 24148 31910 24160
rect 32490 24148 32496 24160
rect 32548 24148 32554 24200
rect 33318 24148 33324 24200
rect 33376 24148 33382 24200
rect 34054 24148 34060 24200
rect 34112 24148 34118 24200
rect 34514 24148 34520 24200
rect 34572 24188 34578 24200
rect 34992 24197 35020 24228
rect 37001 24225 37013 24228
rect 37047 24225 37059 24259
rect 37001 24219 37059 24225
rect 39574 24216 39580 24268
rect 39632 24256 39638 24268
rect 40037 24259 40095 24265
rect 40037 24256 40049 24259
rect 39632 24228 40049 24256
rect 39632 24216 39638 24228
rect 40037 24225 40049 24228
rect 40083 24225 40095 24259
rect 40037 24219 40095 24225
rect 40310 24216 40316 24268
rect 40368 24216 40374 24268
rect 34977 24191 35035 24197
rect 34977 24188 34989 24191
rect 34572 24160 34989 24188
rect 34572 24148 34578 24160
rect 34977 24157 34989 24160
rect 35023 24157 35035 24191
rect 34977 24151 35035 24157
rect 35066 24148 35072 24200
rect 35124 24188 35130 24200
rect 35713 24191 35771 24197
rect 35713 24188 35725 24191
rect 35124 24160 35725 24188
rect 35124 24148 35130 24160
rect 35713 24157 35725 24160
rect 35759 24157 35771 24191
rect 35713 24151 35771 24157
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24188 36599 24191
rect 36814 24188 36820 24200
rect 36587 24160 36820 24188
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 30926 24120 30932 24132
rect 26752 24092 30932 24120
rect 26752 24080 26758 24092
rect 30926 24080 30932 24092
rect 30984 24080 30990 24132
rect 25087 24024 25728 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25774 24012 25780 24064
rect 25832 24012 25838 24064
rect 26142 24012 26148 24064
rect 26200 24012 26206 24064
rect 27154 24012 27160 24064
rect 27212 24012 27218 24064
rect 27246 24012 27252 24064
rect 27304 24052 27310 24064
rect 27525 24055 27583 24061
rect 27525 24052 27537 24055
rect 27304 24024 27537 24052
rect 27304 24012 27310 24024
rect 27525 24021 27537 24024
rect 27571 24021 27583 24055
rect 27525 24015 27583 24021
rect 28350 24012 28356 24064
rect 28408 24012 28414 24064
rect 29546 24012 29552 24064
rect 29604 24052 29610 24064
rect 30837 24055 30895 24061
rect 30837 24052 30849 24055
rect 29604 24024 30849 24052
rect 29604 24012 29610 24024
rect 30837 24021 30849 24024
rect 30883 24021 30895 24055
rect 30837 24015 30895 24021
rect 31386 24012 31392 24064
rect 31444 24052 31450 24064
rect 31757 24055 31815 24061
rect 31757 24052 31769 24055
rect 31444 24024 31769 24052
rect 31444 24012 31450 24024
rect 31757 24021 31769 24024
rect 31803 24021 31815 24055
rect 31757 24015 31815 24021
rect 31846 24012 31852 24064
rect 31904 24052 31910 24064
rect 32309 24055 32367 24061
rect 32309 24052 32321 24055
rect 31904 24024 32321 24052
rect 31904 24012 31910 24024
rect 32309 24021 32321 24024
rect 32355 24021 32367 24055
rect 32309 24015 32367 24021
rect 34606 24012 34612 24064
rect 34664 24052 34670 24064
rect 35069 24055 35127 24061
rect 35069 24052 35081 24055
rect 34664 24024 35081 24052
rect 34664 24012 34670 24024
rect 35069 24021 35081 24024
rect 35115 24021 35127 24055
rect 35728 24052 35756 24151
rect 36814 24148 36820 24160
rect 36872 24148 36878 24200
rect 37274 24148 37280 24200
rect 37332 24188 37338 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 37332 24160 37657 24188
rect 37332 24148 37338 24160
rect 37645 24157 37657 24160
rect 37691 24157 37703 24191
rect 37645 24151 37703 24157
rect 38470 24148 38476 24200
rect 38528 24148 38534 24200
rect 39206 24148 39212 24200
rect 39264 24148 39270 24200
rect 40586 24148 40592 24200
rect 40644 24188 40650 24200
rect 41509 24191 41567 24197
rect 41509 24188 41521 24191
rect 40644 24160 41521 24188
rect 40644 24148 40650 24160
rect 41509 24157 41521 24160
rect 41555 24188 41567 24191
rect 41785 24191 41843 24197
rect 41785 24188 41797 24191
rect 41555 24160 41797 24188
rect 41555 24157 41567 24160
rect 41509 24151 41567 24157
rect 41785 24157 41797 24160
rect 41831 24157 41843 24191
rect 42168 24188 42196 24355
rect 44726 24352 44732 24404
rect 44784 24352 44790 24404
rect 42613 24191 42671 24197
rect 42613 24188 42625 24191
rect 42168 24160 42625 24188
rect 41785 24151 41843 24157
rect 42613 24157 42625 24160
rect 42659 24157 42671 24191
rect 42613 24151 42671 24157
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44784 24160 45201 24188
rect 44784 24148 44790 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45278 24148 45284 24200
rect 45336 24188 45342 24200
rect 45336 24160 45508 24188
rect 45336 24148 45342 24160
rect 35894 24080 35900 24132
rect 35952 24080 35958 24132
rect 37921 24123 37979 24129
rect 37921 24120 37933 24123
rect 36004 24092 37933 24120
rect 36004 24052 36032 24092
rect 37921 24089 37933 24092
rect 37967 24089 37979 24123
rect 37921 24083 37979 24089
rect 40034 24080 40040 24132
rect 40092 24120 40098 24132
rect 45480 24120 45508 24160
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45612 24160 45937 24188
rect 45612 24148 45618 24160
rect 45925 24157 45937 24160
rect 45971 24157 45983 24191
rect 45925 24151 45983 24157
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46661 24191 46719 24197
rect 46661 24188 46673 24191
rect 46072 24160 46673 24188
rect 46072 24148 46078 24160
rect 46661 24157 46673 24160
rect 46707 24188 46719 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 46707 24160 47225 24188
rect 46707 24157 46719 24160
rect 46661 24151 46719 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 47946 24148 47952 24200
rect 48004 24188 48010 24200
rect 48501 24191 48559 24197
rect 48501 24188 48513 24191
rect 48004 24160 48513 24188
rect 48004 24148 48010 24160
rect 48501 24157 48513 24160
rect 48547 24188 48559 24191
rect 49053 24191 49111 24197
rect 49053 24188 49065 24191
rect 48547 24160 49065 24188
rect 48547 24157 48559 24160
rect 48501 24151 48559 24157
rect 49053 24157 49065 24160
rect 49099 24157 49111 24191
rect 49053 24151 49111 24157
rect 40092 24092 43944 24120
rect 45480 24092 47992 24120
rect 40092 24080 40098 24092
rect 35728 24024 36032 24052
rect 35069 24015 35127 24021
rect 36170 24012 36176 24064
rect 36228 24052 36234 24064
rect 36357 24055 36415 24061
rect 36357 24052 36369 24055
rect 36228 24024 36369 24052
rect 36228 24012 36234 24024
rect 36357 24021 36369 24024
rect 36403 24021 36415 24055
rect 36357 24015 36415 24021
rect 37458 24012 37464 24064
rect 37516 24012 37522 24064
rect 39298 24012 39304 24064
rect 39356 24012 39362 24064
rect 41322 24012 41328 24064
rect 41380 24012 41386 24064
rect 43916 24061 43944 24092
rect 43901 24055 43959 24061
rect 43901 24021 43913 24055
rect 43947 24021 43959 24055
rect 43901 24015 43959 24021
rect 43990 24012 43996 24064
rect 44048 24052 44054 24064
rect 45373 24055 45431 24061
rect 45373 24052 45385 24055
rect 44048 24024 45385 24052
rect 44048 24012 44054 24024
rect 45373 24021 45385 24024
rect 45419 24021 45431 24055
rect 45373 24015 45431 24021
rect 45462 24012 45468 24064
rect 45520 24052 45526 24064
rect 46109 24055 46167 24061
rect 46109 24052 46121 24055
rect 45520 24024 46121 24052
rect 45520 24012 45526 24024
rect 46109 24021 46121 24024
rect 46155 24021 46167 24055
rect 46109 24015 46167 24021
rect 46842 24012 46848 24064
rect 46900 24012 46906 24064
rect 47964 24061 47992 24092
rect 47949 24055 48007 24061
rect 47949 24021 47961 24055
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 48682 24012 48688 24064
rect 48740 24012 48746 24064
rect 49510 24012 49516 24064
rect 49568 24012 49574 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 4982 23848 4988 23860
rect 3568 23820 4988 23848
rect 3568 23808 3574 23820
rect 4982 23808 4988 23820
rect 5040 23808 5046 23860
rect 7024 23820 8064 23848
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4154 23780 4160 23792
rect 4019 23752 4160 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23712 2191 23715
rect 2590 23712 2596 23724
rect 2179 23684 2596 23712
rect 2179 23681 2191 23684
rect 2133 23675 2191 23681
rect 2590 23672 2596 23684
rect 2648 23672 2654 23724
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3786 23712 3792 23724
rect 3007 23684 3792 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 7024 23712 7052 23820
rect 7193 23783 7251 23789
rect 7193 23749 7205 23783
rect 7239 23780 7251 23783
rect 7282 23780 7288 23792
rect 7239 23752 7288 23780
rect 7239 23749 7251 23752
rect 7193 23743 7251 23749
rect 7282 23740 7288 23752
rect 7340 23740 7346 23792
rect 4847 23684 7052 23712
rect 7101 23715 7159 23721
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 7101 23681 7113 23715
rect 7147 23681 7159 23715
rect 7101 23675 7159 23681
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6914 23644 6920 23656
rect 5552 23616 6920 23644
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 5552 23576 5580 23616
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 4120 23548 5580 23576
rect 4120 23536 4126 23548
rect 5902 23536 5908 23588
rect 5960 23576 5966 23588
rect 6549 23579 6607 23585
rect 6549 23576 6561 23579
rect 5960 23548 6561 23576
rect 5960 23536 5966 23548
rect 6549 23545 6561 23548
rect 6595 23576 6607 23579
rect 7116 23576 7144 23675
rect 7377 23647 7435 23653
rect 7377 23613 7389 23647
rect 7423 23644 7435 23647
rect 7558 23644 7564 23656
rect 7423 23616 7564 23644
rect 7423 23613 7435 23616
rect 7377 23607 7435 23613
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 8036 23644 8064 23820
rect 12342 23808 12348 23860
rect 12400 23808 12406 23860
rect 17954 23808 17960 23860
rect 18012 23848 18018 23860
rect 21085 23851 21143 23857
rect 21085 23848 21097 23851
rect 18012 23820 21097 23848
rect 18012 23808 18018 23820
rect 21085 23817 21097 23820
rect 21131 23817 21143 23851
rect 21085 23811 21143 23817
rect 21174 23808 21180 23860
rect 21232 23848 21238 23860
rect 24213 23851 24271 23857
rect 21232 23820 24164 23848
rect 21232 23808 21238 23820
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9950 23780 9956 23792
rect 9171 23752 9956 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 12526 23780 12532 23792
rect 11011 23752 12532 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 14185 23783 14243 23789
rect 14185 23749 14197 23783
rect 14231 23780 14243 23783
rect 15746 23780 15752 23792
rect 14231 23752 15752 23780
rect 14231 23749 14243 23752
rect 14185 23743 14243 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 18322 23780 18328 23792
rect 16163 23752 18328 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 18969 23783 19027 23789
rect 18969 23749 18981 23783
rect 19015 23780 19027 23783
rect 19058 23780 19064 23792
rect 19015 23752 19064 23780
rect 19015 23749 19027 23752
rect 18969 23743 19027 23749
rect 19058 23740 19064 23752
rect 19116 23740 19122 23792
rect 20714 23780 20720 23792
rect 20194 23752 20720 23780
rect 20714 23740 20720 23752
rect 20772 23780 20778 23792
rect 21545 23783 21603 23789
rect 21545 23780 21557 23783
rect 20772 23752 21557 23780
rect 20772 23740 20778 23752
rect 21545 23749 21557 23752
rect 21591 23780 21603 23783
rect 22738 23780 22744 23792
rect 21591 23752 22744 23780
rect 21591 23749 21603 23752
rect 21545 23743 21603 23749
rect 22738 23740 22744 23752
rect 22796 23740 22802 23792
rect 24136 23780 24164 23820
rect 24213 23817 24225 23851
rect 24259 23848 24271 23851
rect 24946 23848 24952 23860
rect 24259 23820 24952 23848
rect 24259 23817 24271 23820
rect 24213 23811 24271 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 27154 23848 27160 23860
rect 25056 23820 27160 23848
rect 25056 23780 25084 23820
rect 27154 23808 27160 23820
rect 27212 23808 27218 23860
rect 27706 23808 27712 23860
rect 27764 23848 27770 23860
rect 27764 23820 29684 23848
rect 27764 23808 27770 23820
rect 24136 23752 25084 23780
rect 25590 23740 25596 23792
rect 25648 23740 25654 23792
rect 28166 23740 28172 23792
rect 28224 23740 28230 23792
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23712 8171 23715
rect 8754 23712 8760 23724
rect 8159 23684 8760 23712
rect 8159 23681 8171 23684
rect 8113 23675 8171 23681
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 9858 23672 9864 23724
rect 9916 23672 9922 23724
rect 11793 23715 11851 23721
rect 11793 23681 11805 23715
rect 11839 23712 11851 23715
rect 12250 23712 12256 23724
rect 11839 23684 12256 23712
rect 11839 23681 11851 23684
rect 11793 23675 11851 23681
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 13081 23715 13139 23721
rect 13081 23712 13093 23715
rect 12676 23684 13093 23712
rect 12676 23672 12682 23684
rect 13081 23681 13093 23684
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 14274 23672 14280 23724
rect 14332 23712 14338 23724
rect 14921 23715 14979 23721
rect 14921 23712 14933 23715
rect 14332 23684 14933 23712
rect 14332 23672 14338 23684
rect 14921 23681 14933 23684
rect 14967 23681 14979 23715
rect 14921 23675 14979 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 18138 23712 18144 23724
rect 17083 23684 18144 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18690 23672 18696 23724
rect 18748 23672 18754 23724
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20180 23684 21005 23712
rect 12529 23647 12587 23653
rect 8036 23616 12434 23644
rect 6595 23548 7144 23576
rect 6595 23545 6607 23548
rect 6549 23539 6607 23545
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 2225 23511 2283 23517
rect 2225 23508 2237 23511
rect 1820 23480 2237 23508
rect 1820 23468 1826 23480
rect 2225 23477 2237 23480
rect 2271 23477 2283 23511
rect 2225 23471 2283 23477
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 5258 23508 5264 23520
rect 2832 23480 5264 23508
rect 2832 23468 2838 23480
rect 5258 23468 5264 23480
rect 5316 23468 5322 23520
rect 6178 23468 6184 23520
rect 6236 23508 6242 23520
rect 6365 23511 6423 23517
rect 6365 23508 6377 23511
rect 6236 23480 6377 23508
rect 6236 23468 6242 23480
rect 6365 23477 6377 23480
rect 6411 23477 6423 23511
rect 6365 23471 6423 23477
rect 6730 23468 6736 23520
rect 6788 23468 6794 23520
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 7742 23508 7748 23520
rect 6972 23480 7748 23508
rect 6972 23468 6978 23480
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 11514 23468 11520 23520
rect 11572 23468 11578 23520
rect 11882 23468 11888 23520
rect 11940 23468 11946 23520
rect 12406 23508 12434 23616
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 16942 23644 16948 23656
rect 12575 23616 16948 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 17862 23604 17868 23656
rect 17920 23604 17926 23656
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 20180 23644 20208 23684
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 29546 23672 29552 23724
rect 29604 23672 29610 23724
rect 29656 23712 29684 23820
rect 30926 23808 30932 23860
rect 30984 23808 30990 23860
rect 31110 23808 31116 23860
rect 31168 23848 31174 23860
rect 31297 23851 31355 23857
rect 31297 23848 31309 23851
rect 31168 23820 31309 23848
rect 31168 23808 31174 23820
rect 31297 23817 31309 23820
rect 31343 23817 31355 23851
rect 31297 23811 31355 23817
rect 32858 23808 32864 23860
rect 32916 23848 32922 23860
rect 32953 23851 33011 23857
rect 32953 23848 32965 23851
rect 32916 23820 32965 23848
rect 32916 23808 32922 23820
rect 32953 23817 32965 23820
rect 32999 23817 33011 23851
rect 32953 23811 33011 23817
rect 33594 23808 33600 23860
rect 33652 23848 33658 23860
rect 34057 23851 34115 23857
rect 34057 23848 34069 23851
rect 33652 23820 34069 23848
rect 33652 23808 33658 23820
rect 34057 23817 34069 23820
rect 34103 23817 34115 23851
rect 34057 23811 34115 23817
rect 34790 23808 34796 23860
rect 34848 23808 34854 23860
rect 34974 23808 34980 23860
rect 35032 23848 35038 23860
rect 37458 23848 37464 23860
rect 35032 23820 37464 23848
rect 35032 23808 35038 23820
rect 37458 23808 37464 23820
rect 37516 23808 37522 23860
rect 38470 23808 38476 23860
rect 38528 23808 38534 23860
rect 39025 23851 39083 23857
rect 39025 23817 39037 23851
rect 39071 23848 39083 23851
rect 39206 23848 39212 23860
rect 39071 23820 39212 23848
rect 39071 23817 39083 23820
rect 39025 23811 39083 23817
rect 39206 23808 39212 23820
rect 39264 23808 39270 23860
rect 39574 23808 39580 23860
rect 39632 23848 39638 23860
rect 39853 23851 39911 23857
rect 39853 23848 39865 23851
rect 39632 23820 39865 23848
rect 39632 23808 39638 23820
rect 39853 23817 39865 23820
rect 39899 23817 39911 23851
rect 39853 23811 39911 23817
rect 43257 23851 43315 23857
rect 43257 23817 43269 23851
rect 43303 23848 43315 23851
rect 43438 23848 43444 23860
rect 43303 23820 43444 23848
rect 43303 23817 43315 23820
rect 43257 23811 43315 23817
rect 43438 23808 43444 23820
rect 43496 23808 43502 23860
rect 45554 23808 45560 23860
rect 45612 23848 45618 23860
rect 45741 23851 45799 23857
rect 45741 23848 45753 23851
rect 45612 23820 45753 23848
rect 45612 23808 45618 23820
rect 45741 23817 45753 23820
rect 45787 23817 45799 23851
rect 45741 23811 45799 23817
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 47360 23820 47593 23848
rect 47360 23808 47366 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 30098 23740 30104 23792
rect 30156 23780 30162 23792
rect 33413 23783 33471 23789
rect 33413 23780 33425 23783
rect 30156 23752 33425 23780
rect 30156 23740 30162 23752
rect 33413 23749 33425 23752
rect 33459 23749 33471 23783
rect 35437 23783 35495 23789
rect 35437 23780 35449 23783
rect 33413 23743 33471 23749
rect 33520 23752 35449 23780
rect 29656 23684 31064 23712
rect 19392 23616 20208 23644
rect 22005 23647 22063 23653
rect 19392 23604 19398 23616
rect 22005 23613 22017 23647
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22020 23576 22048 23607
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 23290 23604 23296 23656
rect 23348 23644 23354 23656
rect 24857 23647 24915 23653
rect 24857 23644 24869 23647
rect 23348 23616 24869 23644
rect 23348 23604 23354 23616
rect 24857 23613 24869 23616
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 20088 23548 22048 23576
rect 23753 23579 23811 23585
rect 20088 23520 20116 23548
rect 23753 23545 23765 23579
rect 23799 23576 23811 23579
rect 24394 23576 24400 23588
rect 23799 23548 24400 23576
rect 23799 23545 23811 23548
rect 23753 23539 23811 23545
rect 24394 23536 24400 23548
rect 24452 23536 24458 23588
rect 15102 23508 15108 23520
rect 12406 23480 15108 23508
rect 15102 23468 15108 23480
rect 15160 23468 15166 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 20070 23508 20076 23520
rect 18748 23480 20076 23508
rect 18748 23468 18754 23480
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20441 23511 20499 23517
rect 20441 23477 20453 23511
rect 20487 23508 20499 23511
rect 20530 23508 20536 23520
rect 20487 23480 20536 23508
rect 20487 23477 20499 23480
rect 20441 23471 20499 23477
rect 20530 23468 20536 23480
rect 20588 23468 20594 23520
rect 23842 23468 23848 23520
rect 23900 23508 23906 23520
rect 24578 23508 24584 23520
rect 23900 23480 24584 23508
rect 23900 23468 23906 23480
rect 24578 23468 24584 23480
rect 24636 23468 24642 23520
rect 24872 23508 24900 23607
rect 25130 23604 25136 23656
rect 25188 23604 25194 23656
rect 27154 23644 27160 23656
rect 26160 23616 27160 23644
rect 25682 23508 25688 23520
rect 24872 23480 25688 23508
rect 25682 23468 25688 23480
rect 25740 23508 25746 23520
rect 26160 23508 26188 23616
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 27433 23647 27491 23653
rect 27433 23644 27445 23647
rect 27264 23616 27445 23644
rect 27264 23576 27292 23616
rect 27433 23613 27445 23616
rect 27479 23613 27491 23647
rect 27433 23607 27491 23613
rect 27522 23604 27528 23656
rect 27580 23644 27586 23656
rect 29564 23644 29592 23672
rect 27580 23616 29592 23644
rect 30653 23647 30711 23653
rect 27580 23604 27586 23616
rect 30653 23613 30665 23647
rect 30699 23644 30711 23647
rect 30926 23644 30932 23656
rect 30699 23616 30932 23644
rect 30699 23613 30711 23616
rect 30653 23607 30711 23613
rect 30926 23604 30932 23616
rect 30984 23604 30990 23656
rect 31036 23644 31064 23684
rect 31202 23672 31208 23724
rect 31260 23712 31266 23724
rect 31481 23715 31539 23721
rect 31481 23712 31493 23715
rect 31260 23684 31493 23712
rect 31260 23672 31266 23684
rect 31481 23681 31493 23684
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 32582 23672 32588 23724
rect 32640 23712 32646 23724
rect 33520 23712 33548 23752
rect 35437 23749 35449 23752
rect 35483 23749 35495 23783
rect 35437 23743 35495 23749
rect 35618 23740 35624 23792
rect 35676 23740 35682 23792
rect 32640 23684 33548 23712
rect 33965 23715 34023 23721
rect 32640 23672 32646 23684
rect 33965 23681 33977 23715
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 34701 23715 34759 23721
rect 34701 23681 34713 23715
rect 34747 23712 34759 23715
rect 34882 23712 34888 23724
rect 34747 23684 34888 23712
rect 34747 23681 34759 23684
rect 34701 23675 34759 23681
rect 31846 23644 31852 23656
rect 31036 23616 31852 23644
rect 31846 23604 31852 23616
rect 31904 23604 31910 23656
rect 32309 23647 32367 23653
rect 32309 23613 32321 23647
rect 32355 23613 32367 23647
rect 32309 23607 32367 23613
rect 26620 23548 27292 23576
rect 25740 23480 26188 23508
rect 25740 23468 25746 23480
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 26620 23517 26648 23548
rect 28442 23536 28448 23588
rect 28500 23576 28506 23588
rect 29365 23579 29423 23585
rect 29365 23576 29377 23579
rect 28500 23548 29377 23576
rect 28500 23536 28506 23548
rect 29365 23545 29377 23548
rect 29411 23545 29423 23579
rect 31757 23579 31815 23585
rect 31757 23576 31769 23579
rect 29365 23539 29423 23545
rect 29472 23548 31769 23576
rect 26605 23511 26663 23517
rect 26605 23508 26617 23511
rect 26292 23480 26617 23508
rect 26292 23468 26298 23480
rect 26605 23477 26617 23480
rect 26651 23477 26663 23511
rect 26605 23471 26663 23477
rect 28718 23468 28724 23520
rect 28776 23508 28782 23520
rect 28905 23511 28963 23517
rect 28905 23508 28917 23511
rect 28776 23480 28917 23508
rect 28776 23468 28782 23480
rect 28905 23477 28917 23480
rect 28951 23477 28963 23511
rect 28905 23471 28963 23477
rect 29178 23468 29184 23520
rect 29236 23508 29242 23520
rect 29472 23508 29500 23548
rect 31757 23545 31769 23548
rect 31803 23545 31815 23579
rect 31757 23539 31815 23545
rect 32122 23536 32128 23588
rect 32180 23576 32186 23588
rect 32324 23576 32352 23607
rect 32398 23604 32404 23656
rect 32456 23644 32462 23656
rect 33980 23644 34008 23675
rect 34882 23672 34888 23684
rect 34940 23672 34946 23724
rect 36262 23672 36268 23724
rect 36320 23672 36326 23724
rect 36354 23672 36360 23724
rect 36412 23712 36418 23724
rect 36909 23715 36967 23721
rect 36909 23712 36921 23715
rect 36412 23684 36921 23712
rect 36412 23672 36418 23684
rect 36909 23681 36921 23684
rect 36955 23712 36967 23715
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 36955 23684 37289 23712
rect 36955 23681 36967 23684
rect 36909 23675 36967 23681
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 37642 23672 37648 23724
rect 37700 23712 37706 23724
rect 37921 23715 37979 23721
rect 37921 23712 37933 23715
rect 37700 23684 37933 23712
rect 37700 23672 37706 23684
rect 37921 23681 37933 23684
rect 37967 23712 37979 23715
rect 38197 23715 38255 23721
rect 38197 23712 38209 23715
rect 37967 23684 38209 23712
rect 37967 23681 37979 23684
rect 37921 23675 37979 23681
rect 38197 23681 38209 23684
rect 38243 23681 38255 23715
rect 38197 23675 38255 23681
rect 41138 23672 41144 23724
rect 41196 23712 41202 23724
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 41196 23684 41521 23712
rect 41196 23672 41202 23684
rect 41509 23681 41521 23684
rect 41555 23712 41567 23715
rect 41785 23715 41843 23721
rect 41785 23712 41797 23715
rect 41555 23684 41797 23712
rect 41555 23681 41567 23684
rect 41509 23675 41567 23681
rect 41785 23681 41797 23684
rect 41831 23681 41843 23715
rect 43456 23712 43484 23808
rect 43533 23715 43591 23721
rect 43533 23712 43545 23715
rect 43456 23684 43545 23712
rect 41785 23675 41843 23681
rect 43533 23681 43545 23684
rect 43579 23681 43591 23715
rect 43533 23675 43591 23681
rect 44174 23672 44180 23724
rect 44232 23712 44238 23724
rect 44269 23715 44327 23721
rect 44269 23712 44281 23715
rect 44232 23684 44281 23712
rect 44232 23672 44238 23684
rect 44269 23681 44281 23684
rect 44315 23712 44327 23715
rect 44821 23715 44879 23721
rect 44821 23712 44833 23715
rect 44315 23684 44833 23712
rect 44315 23681 44327 23684
rect 44269 23675 44327 23681
rect 44821 23681 44833 23684
rect 44867 23681 44879 23715
rect 44821 23675 44879 23681
rect 46658 23672 46664 23724
rect 46716 23712 46722 23724
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46716 23684 46765 23712
rect 46716 23672 46722 23684
rect 46753 23681 46765 23684
rect 46799 23712 46811 23715
rect 47305 23715 47363 23721
rect 47305 23712 47317 23715
rect 46799 23684 47317 23712
rect 46799 23681 46811 23684
rect 46753 23675 46811 23681
rect 47305 23681 47317 23684
rect 47351 23681 47363 23715
rect 47305 23675 47363 23681
rect 48041 23715 48099 23721
rect 48041 23681 48053 23715
rect 48087 23712 48099 23715
rect 48314 23712 48320 23724
rect 48087 23684 48320 23712
rect 48087 23681 48099 23684
rect 48041 23675 48099 23681
rect 48314 23672 48320 23684
rect 48372 23672 48378 23724
rect 49053 23715 49111 23721
rect 49053 23681 49065 23715
rect 49099 23712 49111 23715
rect 49510 23712 49516 23724
rect 49099 23684 49516 23712
rect 49099 23681 49111 23684
rect 49053 23675 49111 23681
rect 49510 23672 49516 23684
rect 49568 23672 49574 23724
rect 32456 23616 34008 23644
rect 32456 23604 32462 23616
rect 34606 23604 34612 23656
rect 34664 23644 34670 23656
rect 34664 23616 41368 23644
rect 34664 23604 34670 23616
rect 32180 23548 32352 23576
rect 32180 23536 32186 23548
rect 34698 23536 34704 23588
rect 34756 23576 34762 23588
rect 41340 23585 41368 23616
rect 41598 23604 41604 23656
rect 41656 23644 41662 23656
rect 45462 23644 45468 23656
rect 41656 23616 45468 23644
rect 41656 23604 41662 23616
rect 45462 23604 45468 23616
rect 45520 23604 45526 23656
rect 37737 23579 37795 23585
rect 37737 23576 37749 23579
rect 34756 23548 37749 23576
rect 34756 23536 34762 23548
rect 37737 23545 37749 23548
rect 37783 23545 37795 23579
rect 37737 23539 37795 23545
rect 41325 23579 41383 23585
rect 41325 23545 41337 23579
rect 41371 23545 41383 23579
rect 41325 23539 41383 23545
rect 29236 23480 29500 23508
rect 29236 23468 29242 23480
rect 29546 23468 29552 23520
rect 29604 23508 29610 23520
rect 30193 23511 30251 23517
rect 30193 23508 30205 23511
rect 29604 23480 30205 23508
rect 29604 23468 29610 23480
rect 30193 23477 30205 23480
rect 30239 23477 30251 23511
rect 30193 23471 30251 23477
rect 30466 23468 30472 23520
rect 30524 23508 30530 23520
rect 30745 23511 30803 23517
rect 30745 23508 30757 23511
rect 30524 23480 30757 23508
rect 30524 23468 30530 23480
rect 30745 23477 30757 23480
rect 30791 23477 30803 23511
rect 30745 23471 30803 23477
rect 36078 23468 36084 23520
rect 36136 23468 36142 23520
rect 36722 23468 36728 23520
rect 36780 23468 36786 23520
rect 41414 23468 41420 23520
rect 41472 23508 41478 23520
rect 43717 23511 43775 23517
rect 43717 23508 43729 23511
rect 41472 23480 43729 23508
rect 41472 23468 41478 23480
rect 43717 23477 43729 23480
rect 43763 23477 43775 23511
rect 43717 23471 43775 23477
rect 44450 23468 44456 23520
rect 44508 23468 44514 23520
rect 46934 23468 46940 23520
rect 46992 23468 46998 23520
rect 48498 23468 48504 23520
rect 48556 23468 48562 23520
rect 49234 23468 49240 23520
rect 49292 23468 49298 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 1912 23276 14473 23304
rect 1912 23264 1918 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 17862 23264 17868 23316
rect 17920 23304 17926 23316
rect 19610 23304 19616 23316
rect 17920 23276 19616 23304
rect 17920 23264 17926 23276
rect 19610 23264 19616 23276
rect 19668 23264 19674 23316
rect 19702 23264 19708 23316
rect 19760 23304 19766 23316
rect 22094 23304 22100 23316
rect 19760 23276 22100 23304
rect 19760 23264 19766 23276
rect 22094 23264 22100 23276
rect 22152 23264 22158 23316
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 24302 23304 24308 23316
rect 22244 23276 24308 23304
rect 22244 23264 22250 23276
rect 24302 23264 24308 23276
rect 24360 23264 24366 23316
rect 24394 23264 24400 23316
rect 24452 23304 24458 23316
rect 27512 23307 27570 23313
rect 24452 23276 26372 23304
rect 24452 23264 24458 23276
rect 4157 23239 4215 23245
rect 4157 23205 4169 23239
rect 4203 23236 4215 23239
rect 5166 23236 5172 23248
rect 4203 23208 5172 23236
rect 4203 23205 4215 23208
rect 4157 23199 4215 23205
rect 5166 23196 5172 23208
rect 5224 23196 5230 23248
rect 13722 23196 13728 23248
rect 13780 23236 13786 23248
rect 16574 23236 16580 23248
rect 13780 23208 16580 23236
rect 13780 23196 13786 23208
rect 16574 23196 16580 23208
rect 16632 23196 16638 23248
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19058 23236 19064 23248
rect 18923 23208 19064 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 22278 23236 22284 23248
rect 19352 23208 20208 23236
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 4338 23168 4344 23180
rect 2924 23140 4344 23168
rect 2924 23128 2930 23140
rect 4338 23128 4344 23140
rect 4396 23128 4402 23180
rect 4798 23128 4804 23180
rect 4856 23128 4862 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 12434 23168 12440 23180
rect 11563 23140 12440 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 16485 23171 16543 23177
rect 16485 23137 16497 23171
rect 16531 23168 16543 23171
rect 17402 23168 17408 23180
rect 16531 23140 17408 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 1946 23100 1952 23112
rect 1811 23072 1952 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 1946 23060 1952 23072
rect 2004 23060 2010 23112
rect 3605 23103 3663 23109
rect 3605 23069 3617 23103
rect 3651 23100 3663 23103
rect 4154 23100 4160 23112
rect 3651 23072 4160 23100
rect 3651 23069 3663 23072
rect 3605 23063 3663 23069
rect 4154 23060 4160 23072
rect 4212 23060 4218 23112
rect 4522 23060 4528 23112
rect 4580 23100 4586 23112
rect 4617 23103 4675 23109
rect 4617 23100 4629 23103
rect 4580 23072 4629 23100
rect 4580 23060 4586 23072
rect 4617 23069 4629 23072
rect 4663 23069 4675 23103
rect 4617 23063 4675 23069
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3970 22992 3976 23044
rect 4028 23032 4034 23044
rect 5368 23032 5396 23063
rect 6270 23060 6276 23112
rect 6328 23100 6334 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 6328 23072 7205 23100
rect 6328 23060 6334 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 8352 23072 9321 23100
rect 8352 23060 8358 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 15470 23060 15476 23112
rect 15528 23060 15534 23112
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16908 23072 17141 23100
rect 16908 23060 16914 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 4028 23004 5396 23032
rect 4028 22992 4034 23004
rect 8478 22992 8484 23044
rect 8536 23032 8542 23044
rect 8536 23004 9536 23032
rect 8536 22992 8542 23004
rect 3694 22924 3700 22976
rect 3752 22964 3758 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 3752 22936 3801 22964
rect 3752 22924 3758 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 4065 22967 4123 22973
rect 4065 22933 4077 22967
rect 4111 22964 4123 22967
rect 4525 22967 4583 22973
rect 4525 22964 4537 22967
rect 4111 22936 4537 22964
rect 4111 22933 4123 22936
rect 4065 22927 4123 22933
rect 4525 22933 4537 22936
rect 4571 22964 4583 22967
rect 4706 22964 4712 22976
rect 4571 22936 4712 22964
rect 4571 22933 4583 22936
rect 4525 22927 4583 22933
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 9030 22924 9036 22976
rect 9088 22924 9094 22976
rect 9508 22964 9536 23004
rect 9582 22992 9588 23044
rect 9640 22992 9646 23044
rect 11146 23032 11152 23044
rect 10810 23004 11152 23032
rect 11146 22992 11152 23004
rect 11204 23032 11210 23044
rect 11514 23032 11520 23044
rect 11204 23004 11520 23032
rect 11204 22992 11210 23004
rect 11514 22992 11520 23004
rect 11572 22992 11578 23044
rect 11793 23035 11851 23041
rect 11793 23001 11805 23035
rect 11839 23001 11851 23035
rect 11793 22995 11851 23001
rect 11057 22967 11115 22973
rect 11057 22964 11069 22967
rect 9508 22936 11069 22964
rect 11057 22933 11069 22936
rect 11103 22964 11115 22967
rect 11808 22964 11836 22995
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 11940 23004 12282 23032
rect 11940 22992 11946 23004
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 13633 23035 13691 23041
rect 13633 23032 13645 23035
rect 13228 23004 13645 23032
rect 13228 22992 13234 23004
rect 13633 23001 13645 23004
rect 13679 23032 13691 23035
rect 13814 23032 13820 23044
rect 13679 23004 13820 23032
rect 13679 23001 13691 23004
rect 13633 22995 13691 23001
rect 13814 22992 13820 23004
rect 13872 22992 13878 23044
rect 14366 22992 14372 23044
rect 14424 22992 14430 23044
rect 16942 22992 16948 23044
rect 17000 23032 17006 23044
rect 17405 23035 17463 23041
rect 17405 23032 17417 23035
rect 17000 23004 17417 23032
rect 17000 22992 17006 23004
rect 17405 23001 17417 23004
rect 17451 23001 17463 23035
rect 17405 22995 17463 23001
rect 11103 22936 11836 22964
rect 13265 22967 13323 22973
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 13265 22933 13277 22967
rect 13311 22964 13323 22967
rect 13446 22964 13452 22976
rect 13311 22936 13452 22964
rect 13311 22933 13323 22936
rect 13265 22927 13323 22933
rect 13446 22924 13452 22936
rect 13504 22924 13510 22976
rect 13832 22964 13860 22992
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 13832 22936 14933 22964
rect 14921 22933 14933 22936
rect 14967 22933 14979 22967
rect 14921 22927 14979 22933
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 19352 22964 19380 23208
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 20180 23168 20208 23208
rect 22066 23208 22284 23236
rect 21821 23171 21879 23177
rect 21821 23168 21833 23171
rect 20180 23140 21833 23168
rect 21821 23137 21833 23140
rect 21867 23168 21879 23171
rect 22066 23168 22094 23208
rect 22278 23196 22284 23208
rect 22336 23196 22342 23248
rect 24412 23236 24440 23264
rect 25777 23239 25835 23245
rect 25777 23236 25789 23239
rect 24228 23208 24440 23236
rect 25424 23208 25789 23236
rect 21867 23140 22094 23168
rect 22557 23171 22615 23177
rect 21867 23137 21879 23140
rect 21821 23131 21879 23137
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 24228 23168 24256 23208
rect 22603 23140 24256 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 24302 23128 24308 23180
rect 24360 23168 24366 23180
rect 25133 23171 25191 23177
rect 25133 23168 25145 23171
rect 24360 23140 25145 23168
rect 24360 23128 24366 23140
rect 25133 23137 25145 23140
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23100 19671 23103
rect 19794 23100 19800 23112
rect 19659 23072 19800 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 19794 23060 19800 23072
rect 19852 23060 19858 23112
rect 22278 23060 22284 23112
rect 22336 23060 22342 23112
rect 24118 23060 24124 23112
rect 24176 23100 24182 23112
rect 25424 23100 25452 23208
rect 25777 23205 25789 23208
rect 25823 23205 25835 23239
rect 25777 23199 25835 23205
rect 26344 23177 26372 23276
rect 27512 23273 27524 23307
rect 27558 23304 27570 23307
rect 28718 23304 28724 23316
rect 27558 23276 28724 23304
rect 27558 23273 27570 23276
rect 27512 23267 27570 23273
rect 28718 23264 28724 23276
rect 28776 23264 28782 23316
rect 28994 23264 29000 23316
rect 29052 23304 29058 23316
rect 29990 23307 30048 23313
rect 29990 23304 30002 23307
rect 29052 23276 30002 23304
rect 29052 23264 29058 23276
rect 29990 23273 30002 23276
rect 30036 23273 30048 23307
rect 29990 23267 30048 23273
rect 31202 23264 31208 23316
rect 31260 23304 31266 23316
rect 31941 23307 31999 23313
rect 31941 23304 31953 23307
rect 31260 23276 31953 23304
rect 31260 23264 31266 23276
rect 31941 23273 31953 23276
rect 31987 23273 31999 23307
rect 31941 23267 31999 23273
rect 32030 23264 32036 23316
rect 32088 23304 32094 23316
rect 32493 23307 32551 23313
rect 32493 23304 32505 23307
rect 32088 23276 32505 23304
rect 32088 23264 32094 23276
rect 32493 23273 32505 23276
rect 32539 23273 32551 23307
rect 32493 23267 32551 23273
rect 32674 23264 32680 23316
rect 32732 23304 32738 23316
rect 36262 23304 36268 23316
rect 32732 23276 36268 23304
rect 32732 23264 32738 23276
rect 36262 23264 36268 23276
rect 36320 23304 36326 23316
rect 36633 23307 36691 23313
rect 36633 23304 36645 23307
rect 36320 23276 36645 23304
rect 36320 23264 36326 23276
rect 36633 23273 36645 23276
rect 36679 23273 36691 23307
rect 36633 23267 36691 23273
rect 36814 23264 36820 23316
rect 36872 23264 36878 23316
rect 37274 23264 37280 23316
rect 37332 23264 37338 23316
rect 26988 23208 27384 23236
rect 26329 23171 26387 23177
rect 26329 23137 26341 23171
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 26988 23100 27016 23208
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 27249 23171 27307 23177
rect 27249 23168 27261 23171
rect 27212 23140 27261 23168
rect 27212 23128 27218 23140
rect 27249 23137 27261 23140
rect 27295 23137 27307 23171
rect 27356 23168 27384 23208
rect 28534 23196 28540 23248
rect 28592 23236 28598 23248
rect 28592 23208 29776 23236
rect 28592 23196 28598 23208
rect 27614 23168 27620 23180
rect 27356 23140 27620 23168
rect 27249 23131 27307 23137
rect 27614 23128 27620 23140
rect 27672 23128 27678 23180
rect 28166 23128 28172 23180
rect 28224 23168 28230 23180
rect 29086 23168 29092 23180
rect 28224 23140 29092 23168
rect 28224 23128 28230 23140
rect 29086 23128 29092 23140
rect 29144 23168 29150 23180
rect 29748 23177 29776 23208
rect 31478 23196 31484 23248
rect 31536 23236 31542 23248
rect 34333 23239 34391 23245
rect 34333 23236 34345 23239
rect 31536 23208 34345 23236
rect 31536 23196 31542 23208
rect 34333 23205 34345 23208
rect 34379 23205 34391 23239
rect 34333 23199 34391 23205
rect 35986 23196 35992 23248
rect 36044 23196 36050 23248
rect 29365 23171 29423 23177
rect 29365 23168 29377 23171
rect 29144 23140 29377 23168
rect 29144 23128 29150 23140
rect 29365 23137 29377 23140
rect 29411 23137 29423 23171
rect 29365 23131 29423 23137
rect 29733 23171 29791 23177
rect 29733 23137 29745 23171
rect 29779 23168 29791 23171
rect 37826 23168 37832 23180
rect 29779 23140 37832 23168
rect 29779 23137 29791 23140
rect 29733 23131 29791 23137
rect 24176 23072 25452 23100
rect 25884 23072 27016 23100
rect 24176 23060 24182 23072
rect 20346 22992 20352 23044
rect 20404 22992 20410 23044
rect 20806 22992 20812 23044
rect 20864 22992 20870 23044
rect 22830 22992 22836 23044
rect 22888 23032 22894 23044
rect 22888 23004 23046 23032
rect 22888 22992 22894 23004
rect 16724 22936 19380 22964
rect 19429 22967 19487 22973
rect 16724 22924 16730 22936
rect 19429 22933 19441 22967
rect 19475 22964 19487 22967
rect 20622 22964 20628 22976
rect 19475 22936 20628 22964
rect 19475 22933 19487 22936
rect 19429 22927 19487 22933
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 22940 22964 22968 23004
rect 24762 22992 24768 23044
rect 24820 23032 24826 23044
rect 25590 23032 25596 23044
rect 24820 23004 25596 23032
rect 24820 22992 24826 23004
rect 25590 22992 25596 23004
rect 25648 22992 25654 23044
rect 23290 22964 23296 22976
rect 22940 22936 23296 22964
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 23382 22924 23388 22976
rect 23440 22964 23446 22976
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23440 22936 24041 22964
rect 23440 22924 23446 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24029 22927 24087 22933
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 24946 22924 24952 22976
rect 25004 22924 25010 22976
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25884 22964 25912 23072
rect 26237 23035 26295 23041
rect 26237 23001 26249 23035
rect 26283 23032 26295 23035
rect 26283 23004 27292 23032
rect 26283 23001 26295 23004
rect 26237 22995 26295 23001
rect 25087 22936 25912 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 26142 22924 26148 22976
rect 26200 22964 26206 22976
rect 26510 22964 26516 22976
rect 26200 22936 26516 22964
rect 26200 22924 26206 22936
rect 26510 22924 26516 22936
rect 26568 22964 26574 22976
rect 26789 22967 26847 22973
rect 26789 22964 26801 22967
rect 26568 22936 26801 22964
rect 26568 22924 26574 22936
rect 26789 22933 26801 22936
rect 26835 22933 26847 22967
rect 27264 22964 27292 23004
rect 28166 22992 28172 23044
rect 28224 22992 28230 23044
rect 29380 23032 29408 23131
rect 37826 23128 37832 23140
rect 37884 23128 37890 23180
rect 33321 23103 33379 23109
rect 33321 23069 33333 23103
rect 33367 23100 33379 23103
rect 33686 23100 33692 23112
rect 33367 23072 33692 23100
rect 33367 23069 33379 23072
rect 33321 23063 33379 23069
rect 33686 23060 33692 23072
rect 33744 23060 33750 23112
rect 33778 23060 33784 23112
rect 33836 23100 33842 23112
rect 34057 23103 34115 23109
rect 34057 23100 34069 23103
rect 33836 23072 34069 23100
rect 33836 23060 33842 23072
rect 34057 23069 34069 23072
rect 34103 23069 34115 23103
rect 34057 23063 34115 23069
rect 34422 23060 34428 23112
rect 34480 23100 34486 23112
rect 35069 23103 35127 23109
rect 35069 23100 35081 23103
rect 34480 23072 35081 23100
rect 34480 23060 34486 23072
rect 35069 23069 35081 23072
rect 35115 23069 35127 23103
rect 35069 23063 35127 23069
rect 35710 23060 35716 23112
rect 35768 23060 35774 23112
rect 35986 23060 35992 23112
rect 36044 23100 36050 23112
rect 36173 23103 36231 23109
rect 36173 23100 36185 23103
rect 36044 23072 36185 23100
rect 36044 23060 36050 23072
rect 36173 23069 36185 23072
rect 36219 23069 36231 23103
rect 36173 23063 36231 23069
rect 48590 23060 48596 23112
rect 48648 23060 48654 23112
rect 49053 23103 49111 23109
rect 49053 23069 49065 23103
rect 49099 23100 49111 23103
rect 49326 23100 49332 23112
rect 49099 23072 49332 23100
rect 49099 23069 49111 23072
rect 49053 23063 49111 23069
rect 49326 23060 49332 23072
rect 49384 23060 49390 23112
rect 30006 23032 30012 23044
rect 29380 23004 30012 23032
rect 30006 22992 30012 23004
rect 30064 23032 30070 23044
rect 30466 23032 30472 23044
rect 30064 23004 30472 23032
rect 30064 22992 30070 23004
rect 30466 22992 30472 23004
rect 30524 22992 30530 23044
rect 31312 23004 31892 23032
rect 28350 22964 28356 22976
rect 27264 22936 28356 22964
rect 26789 22927 26847 22933
rect 28350 22924 28356 22936
rect 28408 22924 28414 22976
rect 29730 22924 29736 22976
rect 29788 22964 29794 22976
rect 31312 22964 31340 23004
rect 29788 22936 31340 22964
rect 29788 22924 29794 22936
rect 31478 22924 31484 22976
rect 31536 22924 31542 22976
rect 31662 22924 31668 22976
rect 31720 22964 31726 22976
rect 31757 22967 31815 22973
rect 31757 22964 31769 22967
rect 31720 22936 31769 22964
rect 31720 22924 31726 22936
rect 31757 22933 31769 22936
rect 31803 22933 31815 22967
rect 31864 22964 31892 23004
rect 32122 22992 32128 23044
rect 32180 23032 32186 23044
rect 32401 23035 32459 23041
rect 32401 23032 32413 23035
rect 32180 23004 32413 23032
rect 32180 22992 32186 23004
rect 32401 23001 32413 23004
rect 32447 23001 32459 23035
rect 32401 22995 32459 23001
rect 33137 23035 33195 23041
rect 33137 23001 33149 23035
rect 33183 23032 33195 23035
rect 33410 23032 33416 23044
rect 33183 23004 33416 23032
rect 33183 23001 33195 23004
rect 33137 22995 33195 23001
rect 33410 22992 33416 23004
rect 33468 22992 33474 23044
rect 33873 23035 33931 23041
rect 33873 23001 33885 23035
rect 33919 23001 33931 23035
rect 33873 22995 33931 23001
rect 33888 22964 33916 22995
rect 31864 22936 33916 22964
rect 31757 22927 31815 22933
rect 34514 22924 34520 22976
rect 34572 22964 34578 22976
rect 34885 22967 34943 22973
rect 34885 22964 34897 22967
rect 34572 22936 34897 22964
rect 34572 22924 34578 22936
rect 34885 22933 34897 22936
rect 34931 22933 34943 22967
rect 34885 22927 34943 22933
rect 35526 22924 35532 22976
rect 35584 22924 35590 22976
rect 48406 22924 48412 22976
rect 48464 22924 48470 22976
rect 48774 22924 48780 22976
rect 48832 22964 48838 22976
rect 49237 22967 49295 22973
rect 49237 22964 49249 22967
rect 48832 22936 49249 22964
rect 48832 22924 48838 22936
rect 49237 22933 49249 22936
rect 49283 22933 49295 22967
rect 49237 22927 49295 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 2222 22720 2228 22772
rect 2280 22760 2286 22772
rect 4430 22760 4436 22772
rect 2280 22732 4436 22760
rect 2280 22720 2286 22732
rect 4430 22720 4436 22732
rect 4488 22720 4494 22772
rect 6914 22760 6920 22772
rect 4540 22732 6920 22760
rect 3694 22652 3700 22704
rect 3752 22692 3758 22704
rect 3752 22664 4016 22692
rect 3752 22652 3758 22664
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 1854 22624 1860 22636
rect 1811 22596 1860 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 3602 22584 3608 22636
rect 3660 22624 3666 22636
rect 3789 22627 3847 22633
rect 3789 22624 3801 22627
rect 3660 22596 3801 22624
rect 3660 22584 3666 22596
rect 3789 22593 3801 22596
rect 3835 22593 3847 22627
rect 3988 22624 4016 22664
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 4540 22692 4568 22732
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 9030 22720 9036 22772
rect 9088 22760 9094 22772
rect 14458 22760 14464 22772
rect 9088 22732 14464 22760
rect 9088 22720 9094 22732
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 14645 22763 14703 22769
rect 14645 22729 14657 22763
rect 14691 22760 14703 22763
rect 19702 22760 19708 22772
rect 14691 22732 19708 22760
rect 14691 22729 14703 22732
rect 14645 22723 14703 22729
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 20346 22720 20352 22772
rect 20404 22760 20410 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 20404 22732 21465 22760
rect 20404 22720 20410 22732
rect 21453 22729 21465 22732
rect 21499 22760 21511 22763
rect 22186 22760 22192 22772
rect 21499 22732 22192 22760
rect 21499 22729 21511 22732
rect 21453 22723 21511 22729
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 22465 22763 22523 22769
rect 22465 22729 22477 22763
rect 22511 22760 22523 22763
rect 23658 22760 23664 22772
rect 22511 22732 23664 22760
rect 22511 22729 22523 22732
rect 22465 22723 22523 22729
rect 23658 22720 23664 22732
rect 23716 22720 23722 22772
rect 23768 22732 24532 22760
rect 4120 22664 4568 22692
rect 4632 22664 4936 22692
rect 4120 22652 4126 22664
rect 4632 22624 4660 22664
rect 3988 22596 4660 22624
rect 4801 22627 4859 22633
rect 3789 22587 3847 22593
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4908 22624 4936 22664
rect 5350 22652 5356 22704
rect 5408 22692 5414 22704
rect 5408 22664 7972 22692
rect 5408 22652 5414 22664
rect 6638 22624 6644 22636
rect 4908 22596 6644 22624
rect 4801 22587 4859 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3418 22516 3424 22568
rect 3476 22556 3482 22568
rect 3881 22559 3939 22565
rect 3881 22556 3893 22559
rect 3476 22528 3893 22556
rect 3476 22516 3482 22528
rect 3881 22525 3893 22528
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4062 22516 4068 22568
rect 4120 22516 4126 22568
rect 2406 22448 2412 22500
rect 2464 22488 2470 22500
rect 3970 22488 3976 22500
rect 2464 22460 3976 22488
rect 2464 22448 2470 22460
rect 3970 22448 3976 22460
rect 4028 22448 4034 22500
rect 4816 22488 4844 22587
rect 6638 22584 6644 22596
rect 6696 22584 6702 22636
rect 6730 22584 6736 22636
rect 6788 22624 6794 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 6788 22596 7113 22624
rect 6788 22584 6794 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7650 22624 7656 22636
rect 7239 22596 7656 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 7944 22633 7972 22664
rect 10686 22652 10692 22704
rect 10744 22652 10750 22704
rect 11790 22652 11796 22704
rect 11848 22652 11854 22704
rect 11882 22652 11888 22704
rect 11940 22692 11946 22704
rect 13170 22692 13176 22704
rect 11940 22664 13176 22692
rect 11940 22652 11946 22664
rect 13170 22652 13176 22664
rect 13228 22652 13234 22704
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 17126 22652 17132 22704
rect 17184 22652 17190 22704
rect 18506 22692 18512 22704
rect 18354 22664 18512 22692
rect 18506 22652 18512 22664
rect 18564 22652 18570 22704
rect 20070 22692 20076 22704
rect 19720 22664 20076 22692
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10134 22624 10140 22636
rect 9999 22596 10140 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22624 15163 22627
rect 16758 22624 16764 22636
rect 15151 22596 16764 22624
rect 15151 22593 15163 22596
rect 15105 22587 15163 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19720 22633 19748 22664
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 20714 22652 20720 22704
rect 20772 22652 20778 22704
rect 23290 22692 23296 22704
rect 23124 22664 23296 22692
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19484 22596 19717 22624
rect 19484 22584 19490 22596
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 22278 22584 22284 22636
rect 22336 22624 22342 22636
rect 23124 22633 23152 22664
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 23382 22652 23388 22704
rect 23440 22652 23446 22704
rect 23474 22652 23480 22704
rect 23532 22692 23538 22704
rect 23768 22692 23796 22732
rect 23532 22664 23874 22692
rect 23532 22652 23538 22664
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 22336 22596 23121 22624
rect 22336 22584 22342 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 24504 22624 24532 22732
rect 24670 22720 24676 22772
rect 24728 22760 24734 22772
rect 25682 22760 25688 22772
rect 24728 22732 25688 22760
rect 24728 22720 24734 22732
rect 25682 22720 25688 22732
rect 25740 22720 25746 22772
rect 25777 22763 25835 22769
rect 25777 22729 25789 22763
rect 25823 22760 25835 22763
rect 28442 22760 28448 22772
rect 25823 22732 28448 22760
rect 25823 22729 25835 22732
rect 25777 22723 25835 22729
rect 28442 22720 28448 22732
rect 28500 22720 28506 22772
rect 31478 22760 31484 22772
rect 28644 22732 31484 22760
rect 25130 22652 25136 22704
rect 25188 22692 25194 22704
rect 27338 22692 27344 22704
rect 25188 22664 27344 22692
rect 25188 22652 25194 22664
rect 27338 22652 27344 22664
rect 27396 22692 27402 22704
rect 28534 22692 28540 22704
rect 27396 22664 27660 22692
rect 27396 22652 27402 22664
rect 24762 22624 24768 22636
rect 24504 22610 24768 22624
rect 24518 22596 24768 22610
rect 23109 22587 23167 22593
rect 24762 22584 24768 22596
rect 24820 22584 24826 22636
rect 24946 22584 24952 22636
rect 25004 22624 25010 22636
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25004 22596 25697 22624
rect 25004 22584 25010 22596
rect 25685 22593 25697 22596
rect 25731 22624 25743 22627
rect 26329 22627 26387 22633
rect 26329 22624 26341 22627
rect 25731 22596 26341 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 26329 22593 26341 22596
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 27430 22584 27436 22636
rect 27488 22624 27494 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 27488 22596 27537 22624
rect 27488 22584 27494 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27632 22624 27660 22664
rect 28368 22664 28540 22692
rect 27632 22596 27752 22624
rect 27525 22587 27583 22593
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 7374 22516 7380 22568
rect 7432 22516 7438 22568
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 12434 22516 12440 22568
rect 12492 22516 12498 22568
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22556 12771 22559
rect 13446 22556 13452 22568
rect 12759 22528 13452 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 13446 22516 13452 22528
rect 13504 22516 13510 22568
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 19981 22559 20039 22565
rect 19981 22556 19993 22559
rect 16960 22528 19993 22556
rect 16114 22488 16120 22500
rect 4816 22460 12434 22488
rect 3421 22423 3479 22429
rect 3421 22389 3433 22423
rect 3467 22420 3479 22423
rect 3694 22420 3700 22432
rect 3467 22392 3700 22420
rect 3467 22389 3479 22392
rect 3421 22383 3479 22389
rect 3694 22380 3700 22392
rect 3752 22380 3758 22432
rect 6362 22380 6368 22432
rect 6420 22380 6426 22432
rect 6454 22380 6460 22432
rect 6512 22420 6518 22432
rect 6733 22423 6791 22429
rect 6733 22420 6745 22423
rect 6512 22392 6745 22420
rect 6512 22380 6518 22392
rect 6733 22389 6745 22392
rect 6779 22389 6791 22423
rect 6733 22383 6791 22389
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 7156 22392 11897 22420
rect 7156 22380 7162 22392
rect 11885 22389 11897 22392
rect 11931 22389 11943 22423
rect 12406 22420 12434 22460
rect 14108 22460 16120 22488
rect 14108 22420 14136 22460
rect 16114 22448 16120 22460
rect 16172 22448 16178 22500
rect 16206 22448 16212 22500
rect 16264 22488 16270 22500
rect 16960 22488 16988 22528
rect 19981 22525 19993 22528
rect 20027 22556 20039 22559
rect 20530 22556 20536 22568
rect 20027 22528 20536 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 20622 22516 20628 22568
rect 20680 22556 20686 22568
rect 23382 22556 23388 22568
rect 20680 22528 23388 22556
rect 20680 22516 20686 22528
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 23934 22516 23940 22568
rect 23992 22556 23998 22568
rect 24857 22559 24915 22565
rect 24857 22556 24869 22559
rect 23992 22528 24869 22556
rect 23992 22516 23998 22528
rect 24857 22525 24869 22528
rect 24903 22556 24915 22559
rect 25869 22559 25927 22565
rect 25869 22556 25881 22559
rect 24903 22528 25881 22556
rect 24903 22525 24915 22528
rect 24857 22519 24915 22525
rect 25869 22525 25881 22528
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 27614 22516 27620 22568
rect 27672 22516 27678 22568
rect 27724 22565 27752 22596
rect 28368 22565 28396 22664
rect 28534 22652 28540 22664
rect 28592 22652 28598 22704
rect 28644 22701 28672 22732
rect 31478 22720 31484 22732
rect 31536 22720 31542 22772
rect 31754 22720 31760 22772
rect 31812 22760 31818 22772
rect 32493 22763 32551 22769
rect 32493 22760 32505 22763
rect 31812 22732 32505 22760
rect 31812 22720 31818 22732
rect 32493 22729 32505 22732
rect 32539 22729 32551 22763
rect 32493 22723 32551 22729
rect 33137 22763 33195 22769
rect 33137 22729 33149 22763
rect 33183 22760 33195 22763
rect 33318 22760 33324 22772
rect 33183 22732 33324 22760
rect 33183 22729 33195 22732
rect 33137 22723 33195 22729
rect 33318 22720 33324 22732
rect 33376 22720 33382 22772
rect 39945 22763 40003 22769
rect 39945 22729 39957 22763
rect 39991 22760 40003 22763
rect 40034 22760 40040 22772
rect 39991 22732 40040 22760
rect 39991 22729 40003 22732
rect 39945 22723 40003 22729
rect 28629 22695 28687 22701
rect 28629 22661 28641 22695
rect 28675 22661 28687 22695
rect 28629 22655 28687 22661
rect 29086 22652 29092 22704
rect 29144 22652 29150 22704
rect 31021 22695 31079 22701
rect 31021 22661 31033 22695
rect 31067 22692 31079 22695
rect 36078 22692 36084 22704
rect 31067 22664 36084 22692
rect 31067 22661 31079 22664
rect 31021 22655 31079 22661
rect 36078 22652 36084 22664
rect 36136 22652 36142 22704
rect 39960 22692 39988 22723
rect 40034 22720 40040 22732
rect 40092 22720 40098 22772
rect 48590 22720 48596 22772
rect 48648 22760 48654 22772
rect 48685 22763 48743 22769
rect 48685 22760 48697 22763
rect 48648 22732 48697 22760
rect 48648 22720 48654 22732
rect 48685 22729 48697 22732
rect 48731 22729 48743 22763
rect 48685 22723 48743 22729
rect 49326 22720 49332 22772
rect 49384 22720 49390 22772
rect 39330 22664 39988 22692
rect 30929 22627 30987 22633
rect 30929 22593 30941 22627
rect 30975 22624 30987 22627
rect 31202 22624 31208 22636
rect 30975 22596 31208 22624
rect 30975 22593 30987 22596
rect 30929 22587 30987 22593
rect 31202 22584 31208 22596
rect 31260 22624 31266 22636
rect 31757 22627 31815 22633
rect 31757 22624 31769 22627
rect 31260 22596 31769 22624
rect 31260 22584 31266 22596
rect 31757 22593 31769 22596
rect 31803 22593 31815 22627
rect 31757 22587 31815 22593
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22624 32459 22627
rect 32858 22624 32864 22636
rect 32447 22596 32864 22624
rect 32447 22593 32459 22596
rect 32401 22587 32459 22593
rect 32858 22584 32864 22596
rect 32916 22584 32922 22636
rect 32950 22584 32956 22636
rect 33008 22624 33014 22636
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 33008 22596 33609 22624
rect 33008 22584 33014 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33870 22584 33876 22636
rect 33928 22584 33934 22636
rect 37826 22584 37832 22636
rect 37884 22584 37890 22636
rect 27709 22559 27767 22565
rect 27709 22525 27721 22559
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 28353 22559 28411 22565
rect 28353 22525 28365 22559
rect 28399 22556 28411 22559
rect 28399 22528 28488 22556
rect 28399 22525 28411 22528
rect 28353 22519 28411 22525
rect 16264 22460 16988 22488
rect 18601 22491 18659 22497
rect 16264 22448 16270 22460
rect 18601 22457 18613 22491
rect 18647 22488 18659 22491
rect 18782 22488 18788 22500
rect 18647 22460 18788 22488
rect 18647 22457 18659 22460
rect 18601 22451 18659 22457
rect 18782 22448 18788 22460
rect 18840 22448 18846 22500
rect 24412 22460 24992 22488
rect 12406 22392 14136 22420
rect 11885 22383 11943 22389
rect 14182 22380 14188 22432
rect 14240 22380 14246 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 18414 22420 18420 22432
rect 16816 22392 18420 22420
rect 16816 22380 16822 22392
rect 18414 22380 18420 22392
rect 18472 22380 18478 22432
rect 19061 22423 19119 22429
rect 19061 22389 19073 22423
rect 19107 22420 19119 22423
rect 19150 22420 19156 22432
rect 19107 22392 19156 22420
rect 19107 22389 19119 22392
rect 19061 22383 19119 22389
rect 19150 22380 19156 22392
rect 19208 22380 19214 22432
rect 21818 22380 21824 22432
rect 21876 22420 21882 22432
rect 22005 22423 22063 22429
rect 22005 22420 22017 22423
rect 21876 22392 22017 22420
rect 21876 22380 21882 22392
rect 22005 22389 22017 22392
rect 22051 22420 22063 22423
rect 22097 22423 22155 22429
rect 22097 22420 22109 22423
rect 22051 22392 22109 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22097 22389 22109 22392
rect 22143 22389 22155 22423
rect 22097 22383 22155 22389
rect 23474 22380 23480 22432
rect 23532 22420 23538 22432
rect 24412 22420 24440 22460
rect 23532 22392 24440 22420
rect 24964 22420 24992 22460
rect 25406 22448 25412 22500
rect 25464 22488 25470 22500
rect 27157 22491 27215 22497
rect 27157 22488 27169 22491
rect 25464 22460 27169 22488
rect 25464 22448 25470 22460
rect 27157 22457 27169 22460
rect 27203 22457 27215 22491
rect 27157 22451 27215 22457
rect 28460 22432 28488 22528
rect 28718 22516 28724 22568
rect 28776 22556 28782 22568
rect 31113 22559 31171 22565
rect 31113 22556 31125 22559
rect 28776 22528 31125 22556
rect 28776 22516 28782 22528
rect 31113 22525 31125 22528
rect 31159 22525 31171 22559
rect 31573 22559 31631 22565
rect 31573 22556 31585 22559
rect 31113 22519 31171 22525
rect 31220 22528 31585 22556
rect 30006 22448 30012 22500
rect 30064 22488 30070 22500
rect 31220 22488 31248 22528
rect 31573 22525 31585 22528
rect 31619 22556 31631 22559
rect 31662 22556 31668 22568
rect 31619 22528 31668 22556
rect 31619 22525 31631 22528
rect 31573 22519 31631 22525
rect 31662 22516 31668 22528
rect 31720 22516 31726 22568
rect 33318 22516 33324 22568
rect 33376 22556 33382 22568
rect 38105 22559 38163 22565
rect 33376 22528 35894 22556
rect 33376 22516 33382 22528
rect 30064 22460 31248 22488
rect 30064 22448 30070 22460
rect 31294 22448 31300 22500
rect 31352 22488 31358 22500
rect 35345 22491 35403 22497
rect 35345 22488 35357 22491
rect 31352 22460 35357 22488
rect 31352 22448 31358 22460
rect 35345 22457 35357 22460
rect 35391 22488 35403 22491
rect 35710 22488 35716 22500
rect 35391 22460 35716 22488
rect 35391 22457 35403 22460
rect 35345 22451 35403 22457
rect 35710 22448 35716 22460
rect 35768 22448 35774 22500
rect 25317 22423 25375 22429
rect 25317 22420 25329 22423
rect 24964 22392 25329 22420
rect 23532 22380 23538 22392
rect 25317 22389 25329 22392
rect 25363 22389 25375 22423
rect 25317 22383 25375 22389
rect 26510 22380 26516 22432
rect 26568 22420 26574 22432
rect 26697 22423 26755 22429
rect 26697 22420 26709 22423
rect 26568 22392 26709 22420
rect 26568 22380 26574 22392
rect 26697 22389 26709 22392
rect 26743 22389 26755 22423
rect 26697 22383 26755 22389
rect 28442 22380 28448 22432
rect 28500 22380 28506 22432
rect 29086 22380 29092 22432
rect 29144 22420 29150 22432
rect 30101 22423 30159 22429
rect 30101 22420 30113 22423
rect 29144 22392 30113 22420
rect 29144 22380 29150 22392
rect 30101 22389 30113 22392
rect 30147 22389 30159 22423
rect 30101 22383 30159 22389
rect 30374 22380 30380 22432
rect 30432 22420 30438 22432
rect 30561 22423 30619 22429
rect 30561 22420 30573 22423
rect 30432 22392 30573 22420
rect 30432 22380 30438 22392
rect 30561 22389 30573 22392
rect 30607 22389 30619 22423
rect 30561 22383 30619 22389
rect 32858 22380 32864 22432
rect 32916 22380 32922 22432
rect 33321 22423 33379 22429
rect 33321 22389 33333 22423
rect 33367 22420 33379 22423
rect 33410 22420 33416 22432
rect 33367 22392 33416 22420
rect 33367 22389 33379 22392
rect 33321 22383 33379 22389
rect 33410 22380 33416 22392
rect 33468 22380 33474 22432
rect 34514 22380 34520 22432
rect 34572 22420 34578 22432
rect 34701 22423 34759 22429
rect 34701 22420 34713 22423
rect 34572 22392 34713 22420
rect 34572 22380 34578 22392
rect 34701 22389 34713 22392
rect 34747 22389 34759 22423
rect 34701 22383 34759 22389
rect 34882 22380 34888 22432
rect 34940 22380 34946 22432
rect 35866 22420 35894 22528
rect 38105 22525 38117 22559
rect 38151 22556 38163 22559
rect 48406 22556 48412 22568
rect 38151 22528 48412 22556
rect 38151 22525 38163 22528
rect 38105 22519 38163 22525
rect 48406 22516 48412 22528
rect 48464 22516 48470 22568
rect 39577 22423 39635 22429
rect 39577 22420 39589 22423
rect 35866 22392 39589 22420
rect 39577 22389 39589 22392
rect 39623 22389 39635 22423
rect 39577 22383 39635 22389
rect 49510 22380 49516 22432
rect 49568 22380 49574 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 1946 22176 1952 22228
rect 2004 22216 2010 22228
rect 2004 22188 13492 22216
rect 2004 22176 2010 22188
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 7098 22148 7104 22160
rect 4028 22120 7104 22148
rect 4028 22108 4034 22120
rect 7098 22108 7104 22120
rect 7156 22108 7162 22160
rect 9674 22148 9680 22160
rect 9646 22108 9680 22148
rect 9732 22148 9738 22160
rect 10229 22151 10287 22157
rect 10229 22148 10241 22151
rect 9732 22120 10241 22148
rect 9732 22108 9738 22120
rect 10229 22117 10241 22120
rect 10275 22117 10287 22151
rect 10229 22111 10287 22117
rect 11974 22108 11980 22160
rect 12032 22148 12038 22160
rect 12526 22148 12532 22160
rect 12032 22120 12532 22148
rect 12032 22108 12038 22120
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3292 22052 4445 22080
rect 3292 22040 3298 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 8846 22080 8852 22092
rect 4433 22043 4491 22049
rect 4724 22052 8852 22080
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 3970 22012 3976 22024
rect 1811 21984 3976 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4724 22012 4752 22052
rect 8846 22040 8852 22052
rect 8904 22040 8910 22092
rect 9214 22040 9220 22092
rect 9272 22080 9278 22092
rect 9646 22080 9674 22108
rect 9272 22052 9674 22080
rect 9953 22083 10011 22089
rect 9272 22040 9278 22052
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 10134 22080 10140 22092
rect 9999 22052 10140 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 11238 22040 11244 22092
rect 11296 22040 11302 22092
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 13464 22080 13492 22188
rect 15010 22176 15016 22228
rect 15068 22216 15074 22228
rect 15068 22188 15700 22216
rect 15068 22176 15074 22188
rect 15672 22089 15700 22188
rect 17126 22176 17132 22228
rect 17184 22216 17190 22228
rect 18877 22219 18935 22225
rect 18877 22216 18889 22219
rect 17184 22188 18889 22216
rect 17184 22176 17190 22188
rect 18877 22185 18889 22188
rect 18923 22185 18935 22219
rect 22189 22219 22247 22225
rect 22189 22216 22201 22219
rect 18877 22179 18935 22185
rect 20180 22188 22201 22216
rect 18506 22108 18512 22160
rect 18564 22148 18570 22160
rect 19058 22148 19064 22160
rect 18564 22120 19064 22148
rect 18564 22108 18570 22120
rect 19058 22108 19064 22120
rect 19116 22108 19122 22160
rect 14553 22083 14611 22089
rect 14553 22080 14565 22083
rect 13464 22052 14565 22080
rect 14553 22049 14565 22052
rect 14599 22049 14611 22083
rect 14553 22043 14611 22049
rect 15657 22083 15715 22089
rect 15657 22049 15669 22083
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 19426 22080 19432 22092
rect 17175 22052 19432 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 4111 21984 4752 22012
rect 6273 22015 6331 22021
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 6273 21981 6285 22015
rect 6319 22012 6331 22015
rect 6546 22012 6552 22024
rect 6319 21984 6552 22012
rect 6319 21981 6331 21984
rect 6273 21975 6331 21981
rect 3605 21947 3663 21953
rect 3605 21913 3617 21947
rect 3651 21944 3663 21947
rect 6288 21944 6316 21975
rect 6546 21972 6552 21984
rect 6604 21972 6610 22024
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 22012 7067 22015
rect 7098 22012 7104 22024
rect 7055 21984 7104 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 8757 22015 8815 22021
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 9490 22012 9496 22024
rect 8803 21984 9496 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 10100 21984 10701 22012
rect 10100 21972 10106 21984
rect 10689 21981 10701 21984
rect 10735 22012 10747 22015
rect 10778 22012 10784 22024
rect 10735 21984 10784 22012
rect 10735 21981 10747 21984
rect 10689 21975 10747 21981
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 12802 22012 12808 22024
rect 12575 21984 12808 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 22012 14427 22015
rect 15010 22012 15016 22024
rect 14415 21984 15016 22012
rect 14415 21981 14427 21984
rect 14369 21975 14427 21981
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 15378 21972 15384 22024
rect 15436 21972 15442 22024
rect 18506 21972 18512 22024
rect 18564 21972 18570 22024
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 20180 22012 20208 22188
rect 22189 22185 22201 22188
rect 22235 22216 22247 22219
rect 25038 22216 25044 22228
rect 22235 22188 25044 22216
rect 22235 22185 22247 22188
rect 22189 22179 22247 22185
rect 25038 22176 25044 22188
rect 25096 22176 25102 22228
rect 25148 22188 25360 22216
rect 20254 22108 20260 22160
rect 20312 22148 20318 22160
rect 24670 22148 24676 22160
rect 20312 22120 20944 22148
rect 20312 22108 20318 22120
rect 20916 22089 20944 22120
rect 23952 22120 24676 22148
rect 23952 22089 23980 22120
rect 24670 22108 24676 22120
rect 24728 22108 24734 22160
rect 25148 22089 25176 22188
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 25133 22083 25191 22089
rect 23983 22052 24017 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 25332 22080 25360 22188
rect 28810 22176 28816 22228
rect 28868 22216 28874 22228
rect 34514 22216 34520 22228
rect 28868 22188 34520 22216
rect 28868 22176 28874 22188
rect 34514 22176 34520 22188
rect 34572 22176 34578 22228
rect 40034 22216 40040 22228
rect 35866 22188 40040 22216
rect 27062 22108 27068 22160
rect 27120 22148 27126 22160
rect 27120 22120 27292 22148
rect 27120 22108 27126 22120
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 25332 22052 26065 22080
rect 25133 22043 25191 22049
rect 26053 22049 26065 22052
rect 26099 22080 26111 22083
rect 26418 22080 26424 22092
rect 26099 22052 26424 22080
rect 26099 22049 26111 22052
rect 26053 22043 26111 22049
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 27264 22080 27292 22120
rect 27338 22108 27344 22160
rect 27396 22148 27402 22160
rect 27525 22151 27583 22157
rect 27525 22148 27537 22151
rect 27396 22120 27537 22148
rect 27396 22108 27402 22120
rect 27525 22117 27537 22120
rect 27571 22117 27583 22151
rect 31478 22148 31484 22160
rect 27525 22111 27583 22117
rect 30760 22120 31484 22148
rect 30760 22089 30788 22120
rect 31478 22108 31484 22120
rect 31536 22108 31542 22160
rect 31662 22108 31668 22160
rect 31720 22148 31726 22160
rect 35866 22148 35894 22188
rect 40034 22176 40040 22188
rect 40092 22176 40098 22228
rect 31720 22120 35894 22148
rect 31720 22108 31726 22120
rect 27985 22083 28043 22089
rect 27985 22080 27997 22083
rect 27264 22052 27997 22080
rect 27985 22049 27997 22052
rect 28031 22049 28043 22083
rect 27985 22043 28043 22049
rect 30745 22083 30803 22089
rect 30745 22049 30757 22083
rect 30791 22080 30803 22083
rect 30791 22052 30825 22080
rect 30791 22049 30803 22052
rect 30745 22043 30803 22049
rect 31570 22040 31576 22092
rect 31628 22040 31634 22092
rect 32490 22040 32496 22092
rect 32548 22080 32554 22092
rect 33689 22083 33747 22089
rect 33689 22080 33701 22083
rect 32548 22052 33701 22080
rect 32548 22040 32554 22052
rect 33689 22049 33701 22052
rect 33735 22049 33747 22083
rect 33689 22043 33747 22049
rect 18932 21984 20208 22012
rect 18932 21972 18938 21984
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 25406 22012 25412 22024
rect 23799 21984 25412 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 25406 21972 25412 21984
rect 25464 21972 25470 22024
rect 25590 21972 25596 22024
rect 25648 22012 25654 22024
rect 25777 22015 25835 22021
rect 25777 22012 25789 22015
rect 25648 21984 25789 22012
rect 25648 21972 25654 21984
rect 25777 21981 25789 21984
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 27856 21984 28825 22012
rect 27856 21972 27862 21984
rect 28813 21981 28825 21984
rect 28859 22012 28871 22015
rect 29273 22015 29331 22021
rect 29273 22012 29285 22015
rect 28859 21984 29285 22012
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 29273 21981 29285 21984
rect 29319 21981 29331 22015
rect 29273 21975 29331 21981
rect 29825 22015 29883 22021
rect 29825 21981 29837 22015
rect 29871 22012 29883 22015
rect 30561 22015 30619 22021
rect 29871 21984 30512 22012
rect 29871 21981 29883 21984
rect 29825 21975 29883 21981
rect 30484 21956 30512 21984
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 30607 21984 32076 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 3651 21916 6316 21944
rect 3651 21913 3663 21916
rect 3605 21907 3663 21913
rect 6822 21904 6828 21956
rect 6880 21944 6886 21956
rect 7837 21947 7895 21953
rect 7837 21944 7849 21947
rect 6880 21916 7849 21944
rect 6880 21904 6886 21916
rect 7837 21913 7849 21916
rect 7883 21913 7895 21947
rect 7837 21907 7895 21913
rect 8573 21947 8631 21953
rect 8573 21913 8585 21947
rect 8619 21944 8631 21947
rect 11790 21944 11796 21956
rect 8619 21916 11796 21944
rect 8619 21913 8631 21916
rect 8573 21907 8631 21913
rect 11790 21904 11796 21916
rect 11848 21904 11854 21956
rect 17405 21947 17463 21953
rect 17405 21913 17417 21947
rect 17451 21944 17463 21947
rect 17494 21944 17500 21956
rect 17451 21916 17500 21944
rect 17451 21913 17463 21916
rect 17405 21907 17463 21913
rect 17494 21904 17500 21916
rect 17552 21904 17558 21956
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21913 19579 21947
rect 19521 21907 19579 21913
rect 3329 21879 3387 21885
rect 3329 21845 3341 21879
rect 3375 21876 3387 21879
rect 3418 21876 3424 21888
rect 3375 21848 3424 21876
rect 3375 21845 3387 21848
rect 3329 21839 3387 21845
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 5810 21836 5816 21888
rect 5868 21836 5874 21888
rect 6086 21836 6092 21888
rect 6144 21836 6150 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 8386 21876 8392 21888
rect 7800 21848 8392 21876
rect 7800 21836 7806 21848
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 8938 21836 8944 21888
rect 8996 21836 9002 21888
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 9398 21876 9404 21888
rect 9355 21848 9404 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 9769 21879 9827 21885
rect 9769 21845 9781 21879
rect 9815 21876 9827 21879
rect 11422 21876 11428 21888
rect 9815 21848 11428 21876
rect 9815 21845 9827 21848
rect 9769 21839 9827 21845
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 11514 21836 11520 21888
rect 11572 21876 11578 21888
rect 14921 21879 14979 21885
rect 14921 21876 14933 21879
rect 11572 21848 14933 21876
rect 11572 21836 11578 21848
rect 14921 21845 14933 21848
rect 14967 21876 14979 21879
rect 19536 21876 19564 21907
rect 19978 21904 19984 21956
rect 20036 21944 20042 21956
rect 21358 21944 21364 21956
rect 20036 21916 21364 21944
rect 20036 21904 20042 21916
rect 21358 21904 21364 21916
rect 21416 21904 21422 21956
rect 22649 21947 22707 21953
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 22695 21916 24961 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 25222 21904 25228 21956
rect 25280 21944 25286 21956
rect 26510 21944 26516 21956
rect 25280 21916 26516 21944
rect 25280 21904 25286 21916
rect 26510 21904 26516 21916
rect 26568 21904 26574 21956
rect 28994 21904 29000 21956
rect 29052 21944 29058 21956
rect 29052 21916 30144 21944
rect 29052 21904 29058 21916
rect 14967 21848 19564 21876
rect 14967 21845 14979 21848
rect 14921 21839 14979 21845
rect 19610 21836 19616 21888
rect 19668 21836 19674 21888
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 21726 21876 21732 21888
rect 20128 21848 21732 21876
rect 20128 21836 20134 21848
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 22094 21836 22100 21888
rect 22152 21836 22158 21888
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 23293 21879 23351 21885
rect 23293 21876 23305 21879
rect 22428 21848 23305 21876
rect 22428 21836 22434 21848
rect 23293 21845 23305 21848
rect 23339 21845 23351 21879
rect 23293 21839 23351 21845
rect 23658 21836 23664 21888
rect 23716 21836 23722 21888
rect 24578 21836 24584 21888
rect 24636 21836 24642 21888
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 27338 21876 27344 21888
rect 25087 21848 27344 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 28350 21836 28356 21888
rect 28408 21876 28414 21888
rect 28534 21876 28540 21888
rect 28408 21848 28540 21876
rect 28408 21836 28414 21848
rect 28534 21836 28540 21848
rect 28592 21836 28598 21888
rect 28626 21836 28632 21888
rect 28684 21836 28690 21888
rect 29178 21836 29184 21888
rect 29236 21876 29242 21888
rect 29549 21879 29607 21885
rect 29549 21876 29561 21879
rect 29236 21848 29561 21876
rect 29236 21836 29242 21848
rect 29549 21845 29561 21848
rect 29595 21876 29607 21879
rect 30006 21876 30012 21888
rect 29595 21848 30012 21876
rect 29595 21845 29607 21848
rect 29549 21839 29607 21845
rect 30006 21836 30012 21848
rect 30064 21836 30070 21888
rect 30116 21885 30144 21916
rect 30466 21904 30472 21956
rect 30524 21944 30530 21956
rect 31294 21944 31300 21956
rect 30524 21916 31300 21944
rect 30524 21904 30530 21916
rect 31294 21904 31300 21916
rect 31352 21904 31358 21956
rect 31389 21947 31447 21953
rect 31389 21913 31401 21947
rect 31435 21944 31447 21947
rect 31849 21947 31907 21953
rect 31849 21944 31861 21947
rect 31435 21916 31861 21944
rect 31435 21913 31447 21916
rect 31389 21907 31447 21913
rect 31849 21913 31861 21916
rect 31895 21913 31907 21947
rect 32048 21944 32076 21984
rect 32122 21972 32128 22024
rect 32180 22012 32186 22024
rect 32585 22015 32643 22021
rect 32585 22012 32597 22015
rect 32180 21984 32597 22012
rect 32180 21972 32186 21984
rect 32585 21981 32597 21984
rect 32631 21981 32643 22015
rect 32585 21975 32643 21981
rect 32766 21972 32772 22024
rect 32824 22012 32830 22024
rect 32861 22015 32919 22021
rect 32861 22012 32873 22015
rect 32824 21984 32873 22012
rect 32824 21972 32830 21984
rect 32861 21981 32873 21984
rect 32907 21981 32919 22015
rect 32861 21975 32919 21981
rect 49053 22015 49111 22021
rect 49053 21981 49065 22015
rect 49099 22012 49111 22015
rect 49510 22012 49516 22024
rect 49099 21984 49516 22012
rect 49099 21981 49111 21984
rect 49053 21975 49111 21981
rect 49510 21972 49516 21984
rect 49568 21972 49574 22024
rect 36170 21944 36176 21956
rect 32048 21916 36176 21944
rect 31849 21907 31907 21913
rect 30101 21879 30159 21885
rect 30101 21845 30113 21879
rect 30147 21845 30159 21879
rect 30101 21839 30159 21845
rect 31018 21836 31024 21888
rect 31076 21876 31082 21888
rect 31404 21876 31432 21907
rect 36170 21904 36176 21916
rect 36228 21904 36234 21956
rect 31076 21848 31432 21876
rect 31076 21836 31082 21848
rect 32030 21836 32036 21888
rect 32088 21876 32094 21888
rect 32125 21879 32183 21885
rect 32125 21876 32137 21879
rect 32088 21848 32137 21876
rect 32088 21836 32094 21848
rect 32125 21845 32137 21848
rect 32171 21845 32183 21879
rect 32125 21839 32183 21845
rect 48314 21836 48320 21888
rect 48372 21876 48378 21888
rect 49237 21879 49295 21885
rect 49237 21876 49249 21879
rect 48372 21848 49249 21876
rect 48372 21836 48378 21848
rect 49237 21845 49249 21848
rect 49283 21845 49295 21879
rect 49237 21839 49295 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 5534 21672 5540 21684
rect 1780 21644 5540 21672
rect 1780 21545 1808 21644
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 9401 21675 9459 21681
rect 7024 21644 9352 21672
rect 4338 21564 4344 21616
rect 4396 21564 4402 21616
rect 5810 21564 5816 21616
rect 5868 21604 5874 21616
rect 7024 21613 7052 21644
rect 7009 21607 7067 21613
rect 7009 21604 7021 21607
rect 5868 21576 7021 21604
rect 5868 21564 5874 21576
rect 7009 21573 7021 21576
rect 7055 21573 7067 21607
rect 7009 21567 7067 21573
rect 7558 21564 7564 21616
rect 7616 21604 7622 21616
rect 7834 21604 7840 21616
rect 7616 21576 7840 21604
rect 7616 21564 7622 21576
rect 7834 21564 7840 21576
rect 7892 21604 7898 21616
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 7892 21576 7941 21604
rect 7892 21564 7898 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 7929 21567 7987 21573
rect 8938 21564 8944 21616
rect 8996 21564 9002 21616
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 2222 21496 2228 21548
rect 2280 21536 2286 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2280 21508 3433 21536
rect 2280 21496 2286 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 1452 21440 2053 21468
rect 1452 21428 1458 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 2041 21431 2099 21437
rect 2746 21440 5733 21468
rect 2130 21360 2136 21412
rect 2188 21400 2194 21412
rect 2746 21400 2774 21440
rect 5721 21437 5733 21440
rect 5767 21437 5779 21471
rect 5721 21431 5779 21437
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6638 21468 6644 21480
rect 5951 21440 6644 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 7642 21471 7700 21477
rect 7642 21468 7654 21471
rect 7576 21440 7654 21468
rect 2188 21372 2774 21400
rect 2188 21360 2194 21372
rect 4890 21360 4896 21412
rect 4948 21400 4954 21412
rect 7193 21403 7251 21409
rect 7193 21400 7205 21403
rect 4948 21372 7205 21400
rect 4948 21360 4954 21372
rect 7193 21369 7205 21372
rect 7239 21369 7251 21403
rect 7193 21363 7251 21369
rect 5261 21335 5319 21341
rect 5261 21301 5273 21335
rect 5307 21332 5319 21335
rect 5534 21332 5540 21344
rect 5307 21304 5540 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 6362 21292 6368 21344
rect 6420 21292 6426 21344
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 7006 21332 7012 21344
rect 6687 21304 7012 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 7576 21332 7604 21440
rect 7642 21437 7654 21440
rect 7688 21437 7700 21471
rect 7642 21431 7700 21437
rect 9324 21400 9352 21644
rect 9401 21641 9413 21675
rect 9447 21641 9459 21675
rect 9401 21635 9459 21641
rect 9416 21604 9444 21635
rect 9490 21632 9496 21684
rect 9548 21672 9554 21684
rect 9766 21672 9772 21684
rect 9548 21644 9772 21672
rect 9548 21632 9554 21644
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 12158 21672 12164 21684
rect 9907 21644 12164 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 14182 21672 14188 21684
rect 13372 21644 14188 21672
rect 9582 21604 9588 21616
rect 9416 21576 9588 21604
rect 9582 21564 9588 21576
rect 9640 21604 9646 21616
rect 9640 21576 12296 21604
rect 9640 21564 9646 21576
rect 9766 21496 9772 21548
rect 9824 21536 9830 21548
rect 10229 21539 10287 21545
rect 10229 21536 10241 21539
rect 9824 21508 10241 21536
rect 9824 21496 9830 21508
rect 10229 21505 10241 21508
rect 10275 21536 10287 21539
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 10275 21508 10701 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10689 21505 10701 21508
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 11146 21496 11152 21548
rect 11204 21536 11210 21548
rect 11241 21539 11299 21545
rect 11241 21536 11253 21539
rect 11204 21508 11253 21536
rect 11204 21496 11210 21508
rect 11241 21505 11253 21508
rect 11287 21505 11299 21539
rect 11241 21499 11299 21505
rect 11974 21496 11980 21548
rect 12032 21536 12038 21548
rect 12161 21539 12219 21545
rect 12161 21536 12173 21539
rect 12032 21508 12173 21536
rect 12032 21496 12038 21508
rect 12161 21505 12173 21508
rect 12207 21505 12219 21539
rect 12268 21536 12296 21576
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 13372 21613 13400 21644
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 15473 21675 15531 21681
rect 15473 21641 15485 21675
rect 15519 21672 15531 21675
rect 15930 21672 15936 21684
rect 15519 21644 15936 21672
rect 15519 21641 15531 21644
rect 15473 21635 15531 21641
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 16025 21675 16083 21681
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 17678 21672 17684 21684
rect 16071 21644 17684 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 17770 21632 17776 21684
rect 17828 21672 17834 21684
rect 20254 21672 20260 21684
rect 17828 21644 20260 21672
rect 17828 21632 17834 21644
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 23474 21672 23480 21684
rect 22511 21644 23480 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 24578 21672 24584 21684
rect 23584 21644 24584 21672
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 12400 21576 13369 21604
rect 12400 21564 12406 21576
rect 13357 21573 13369 21576
rect 13403 21573 13415 21607
rect 13357 21567 13415 21573
rect 13814 21564 13820 21616
rect 13872 21564 13878 21616
rect 15378 21564 15384 21616
rect 15436 21604 15442 21616
rect 18506 21604 18512 21616
rect 15436 21576 18512 21604
rect 15436 21564 15442 21576
rect 18506 21564 18512 21576
rect 18564 21564 18570 21616
rect 20714 21604 20720 21616
rect 20194 21590 20720 21604
rect 20180 21576 20720 21590
rect 12268 21508 12388 21536
rect 12161 21499 12219 21505
rect 9858 21428 9864 21480
rect 9916 21468 9922 21480
rect 10321 21471 10379 21477
rect 10321 21468 10333 21471
rect 9916 21440 10333 21468
rect 9916 21428 9922 21440
rect 10321 21437 10333 21440
rect 10367 21437 10379 21471
rect 10321 21431 10379 21437
rect 10413 21471 10471 21477
rect 10413 21437 10425 21471
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 10965 21471 11023 21477
rect 10965 21437 10977 21471
rect 11011 21468 11023 21471
rect 12250 21468 12256 21480
rect 11011 21440 12256 21468
rect 11011 21437 11023 21440
rect 10965 21431 11023 21437
rect 10226 21400 10232 21412
rect 9324 21372 10232 21400
rect 10226 21360 10232 21372
rect 10284 21360 10290 21412
rect 10428 21400 10456 21431
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12360 21477 12388 21508
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12492 21508 13093 21536
rect 12492 21496 12498 21508
rect 13081 21505 13093 21508
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 15102 21496 15108 21548
rect 15160 21536 15166 21548
rect 16666 21536 16672 21548
rect 15160 21508 16672 21536
rect 15160 21496 15166 21508
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 17034 21496 17040 21548
rect 17092 21496 17098 21548
rect 12345 21471 12403 21477
rect 12345 21437 12357 21471
rect 12391 21437 12403 21471
rect 13446 21468 13452 21480
rect 12345 21431 12403 21437
rect 12452 21440 13452 21468
rect 12452 21400 12480 21440
rect 13446 21428 13452 21440
rect 13504 21468 13510 21480
rect 13504 21440 15700 21468
rect 13504 21428 13510 21440
rect 10428 21372 12480 21400
rect 14458 21360 14464 21412
rect 14516 21400 14522 21412
rect 15197 21403 15255 21409
rect 15197 21400 15209 21403
rect 14516 21372 15209 21400
rect 14516 21360 14522 21372
rect 15197 21369 15209 21372
rect 15243 21400 15255 21403
rect 15286 21400 15292 21412
rect 15243 21372 15292 21400
rect 15243 21369 15255 21372
rect 15197 21363 15255 21369
rect 15286 21360 15292 21372
rect 15344 21360 15350 21412
rect 15562 21360 15568 21412
rect 15620 21360 15626 21412
rect 15672 21400 15700 21440
rect 16206 21428 16212 21480
rect 16264 21428 16270 21480
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21468 18751 21471
rect 18739 21440 18828 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 17678 21400 17684 21412
rect 15672 21372 17684 21400
rect 17678 21360 17684 21372
rect 17736 21360 17742 21412
rect 8294 21332 8300 21344
rect 7576 21304 8300 21332
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 9766 21292 9772 21344
rect 9824 21292 9830 21344
rect 11790 21292 11796 21344
rect 11848 21292 11854 21344
rect 14829 21335 14887 21341
rect 14829 21301 14841 21335
rect 14875 21332 14887 21335
rect 15010 21332 15016 21344
rect 14875 21304 15016 21332
rect 14875 21301 14887 21304
rect 14829 21295 14887 21301
rect 15010 21292 15016 21304
rect 15068 21292 15074 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 18598 21332 18604 21344
rect 15712 21304 18604 21332
rect 15712 21292 15718 21304
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 18800 21332 18828 21440
rect 18966 21428 18972 21480
rect 19024 21428 19030 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 20180 21468 20208 21576
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 23584 21604 23612 21644
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 25961 21675 26019 21681
rect 25961 21641 25973 21675
rect 26007 21672 26019 21675
rect 27062 21672 27068 21684
rect 26007 21644 27068 21672
rect 26007 21641 26019 21644
rect 25961 21635 26019 21641
rect 27062 21632 27068 21644
rect 27120 21632 27126 21684
rect 27249 21675 27307 21681
rect 27249 21641 27261 21675
rect 27295 21672 27307 21675
rect 27338 21672 27344 21684
rect 27295 21644 27344 21672
rect 27295 21641 27307 21644
rect 27249 21635 27307 21641
rect 27338 21632 27344 21644
rect 27396 21632 27402 21684
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 35526 21672 35532 21684
rect 27755 21644 35532 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 35526 21632 35532 21644
rect 35584 21632 35590 21684
rect 36538 21632 36544 21684
rect 36596 21672 36602 21684
rect 46934 21672 46940 21684
rect 36596 21644 46940 21672
rect 36596 21632 36602 21644
rect 46934 21632 46940 21644
rect 46992 21632 46998 21684
rect 23216 21576 23612 21604
rect 23661 21607 23719 21613
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21315 21508 22385 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 23216 21536 23244 21576
rect 23661 21573 23673 21607
rect 23707 21604 23719 21607
rect 23934 21604 23940 21616
rect 23707 21576 23940 21604
rect 23707 21573 23719 21576
rect 23661 21567 23719 21573
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 25130 21564 25136 21616
rect 25188 21604 25194 21616
rect 26053 21607 26111 21613
rect 25188 21576 25544 21604
rect 25188 21564 25194 21576
rect 22373 21499 22431 21505
rect 22480 21508 23244 21536
rect 19116 21440 20208 21468
rect 19116 21428 19122 21440
rect 20346 21428 20352 21480
rect 20404 21468 20410 21480
rect 22480 21468 22508 21508
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23348 21508 23397 21536
rect 23348 21496 23354 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 24762 21496 24768 21548
rect 24820 21536 24826 21548
rect 25222 21536 25228 21548
rect 24820 21508 25228 21536
rect 24820 21496 24826 21508
rect 25222 21496 25228 21508
rect 25280 21496 25286 21548
rect 25516 21536 25544 21576
rect 26053 21573 26065 21607
rect 26099 21604 26111 21607
rect 28994 21604 29000 21616
rect 26099 21576 29000 21604
rect 26099 21573 26111 21576
rect 26053 21567 26111 21573
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 29178 21564 29184 21616
rect 29236 21564 29242 21616
rect 31113 21607 31171 21613
rect 31113 21573 31125 21607
rect 31159 21604 31171 21607
rect 36722 21604 36728 21616
rect 31159 21576 36728 21604
rect 31159 21573 31171 21576
rect 31113 21567 31171 21573
rect 36722 21564 36728 21576
rect 36780 21564 36786 21616
rect 26697 21539 26755 21545
rect 26697 21536 26709 21539
rect 25516 21508 26709 21536
rect 26697 21505 26709 21508
rect 26743 21536 26755 21539
rect 27617 21539 27675 21545
rect 27617 21536 27629 21539
rect 26743 21508 27629 21536
rect 26743 21505 26755 21508
rect 26697 21499 26755 21505
rect 27617 21505 27629 21508
rect 27663 21536 27675 21539
rect 28074 21536 28080 21548
rect 27663 21508 28080 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 28350 21496 28356 21548
rect 28408 21536 28414 21548
rect 28445 21539 28503 21545
rect 28445 21536 28457 21539
rect 28408 21508 28457 21536
rect 28408 21496 28414 21508
rect 28445 21505 28457 21508
rect 28491 21505 28503 21539
rect 28445 21499 28503 21505
rect 30926 21496 30932 21548
rect 30984 21536 30990 21548
rect 31021 21539 31079 21545
rect 31021 21536 31033 21539
rect 30984 21508 31033 21536
rect 30984 21496 30990 21508
rect 31021 21505 31033 21508
rect 31067 21505 31079 21539
rect 31021 21499 31079 21505
rect 31754 21496 31760 21548
rect 31812 21496 31818 21548
rect 32398 21496 32404 21548
rect 32456 21496 32462 21548
rect 47854 21496 47860 21548
rect 47912 21536 47918 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47912 21508 47961 21536
rect 47912 21496 47918 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 20404 21440 22508 21468
rect 22649 21471 22707 21477
rect 20404 21428 20410 21440
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 24670 21468 24676 21480
rect 22695 21440 24676 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 24670 21428 24676 21440
rect 24728 21468 24734 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24728 21440 25145 21468
rect 24728 21428 24734 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21437 26295 21471
rect 26237 21431 26295 21437
rect 20806 21360 20812 21412
rect 20864 21400 20870 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 20864 21372 22017 21400
rect 20864 21360 20870 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 26252 21400 26280 21431
rect 27890 21428 27896 21480
rect 27948 21428 27954 21480
rect 28721 21471 28779 21477
rect 28721 21468 28733 21471
rect 28552 21440 28733 21468
rect 28552 21400 28580 21440
rect 28721 21437 28733 21440
rect 28767 21468 28779 21471
rect 29086 21468 29092 21480
rect 28767 21440 29092 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 29086 21428 29092 21440
rect 29144 21428 29150 21480
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 30208 21440 31217 21468
rect 26252 21372 28580 21400
rect 22005 21363 22063 21369
rect 19426 21332 19432 21344
rect 18800 21304 19432 21332
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 19760 21304 20453 21332
rect 19760 21292 19766 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 20441 21295 20499 21301
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 20993 21335 21051 21341
rect 20993 21332 21005 21335
rect 20772 21304 21005 21332
rect 20772 21292 20778 21304
rect 20993 21301 21005 21304
rect 21039 21332 21051 21335
rect 21818 21332 21824 21344
rect 21039 21304 21824 21332
rect 21039 21301 21051 21304
rect 20993 21295 21051 21301
rect 21818 21292 21824 21304
rect 21876 21332 21882 21344
rect 23017 21335 23075 21341
rect 23017 21332 23029 21335
rect 21876 21304 23029 21332
rect 21876 21292 21882 21304
rect 23017 21301 23029 21304
rect 23063 21301 23075 21335
rect 23017 21295 23075 21301
rect 23474 21292 23480 21344
rect 23532 21332 23538 21344
rect 24210 21332 24216 21344
rect 23532 21304 24216 21332
rect 23532 21292 23538 21304
rect 24210 21292 24216 21304
rect 24268 21292 24274 21344
rect 24302 21292 24308 21344
rect 24360 21332 24366 21344
rect 25593 21335 25651 21341
rect 25593 21332 25605 21335
rect 24360 21304 25605 21332
rect 24360 21292 24366 21304
rect 25593 21301 25605 21304
rect 25639 21301 25651 21335
rect 25593 21295 25651 21301
rect 28902 21292 28908 21344
rect 28960 21332 28966 21344
rect 30208 21341 30236 21440
rect 31205 21437 31217 21440
rect 31251 21437 31263 21471
rect 31205 21431 31263 21437
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 30282 21360 30288 21412
rect 30340 21400 30346 21412
rect 32122 21400 32128 21412
rect 30340 21372 32128 21400
rect 30340 21360 30346 21372
rect 32122 21360 32128 21372
rect 32180 21360 32186 21412
rect 32674 21360 32680 21412
rect 32732 21400 32738 21412
rect 48498 21400 48504 21412
rect 32732 21372 48504 21400
rect 32732 21360 32738 21372
rect 48498 21360 48504 21372
rect 48556 21360 48562 21412
rect 30193 21335 30251 21341
rect 30193 21332 30205 21335
rect 28960 21304 30205 21332
rect 28960 21292 28966 21304
rect 30193 21301 30205 21304
rect 30239 21301 30251 21335
rect 30193 21295 30251 21301
rect 30650 21292 30656 21344
rect 30708 21292 30714 21344
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 31849 21335 31907 21341
rect 31849 21332 31861 21335
rect 30984 21304 31861 21332
rect 30984 21292 30990 21304
rect 31849 21301 31861 21304
rect 31895 21301 31907 21335
rect 31849 21295 31907 21301
rect 32490 21292 32496 21344
rect 32548 21292 32554 21344
rect 47673 21335 47731 21341
rect 47673 21301 47685 21335
rect 47719 21332 47731 21335
rect 47854 21332 47860 21344
rect 47719 21304 47860 21332
rect 47719 21301 47731 21304
rect 47673 21295 47731 21301
rect 47854 21292 47860 21304
rect 47912 21292 47918 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 3476 21100 7328 21128
rect 3476 21088 3482 21100
rect 7300 21060 7328 21100
rect 7374 21088 7380 21140
rect 7432 21128 7438 21140
rect 8570 21128 8576 21140
rect 7432 21100 8576 21128
rect 7432 21088 7438 21100
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 11514 21128 11520 21140
rect 8720 21100 11520 21128
rect 8720 21088 8726 21100
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 13817 21131 13875 21137
rect 13817 21128 13829 21131
rect 12176 21100 13829 21128
rect 7300 21032 8248 21060
rect 3881 20995 3939 21001
rect 3881 20961 3893 20995
rect 3927 20992 3939 20995
rect 3970 20992 3976 21004
rect 3927 20964 3976 20992
rect 3927 20961 3939 20964
rect 3881 20955 3939 20961
rect 3970 20952 3976 20964
rect 4028 20952 4034 21004
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 5721 20995 5779 21001
rect 5721 20961 5733 20995
rect 5767 20992 5779 20995
rect 7374 20992 7380 21004
rect 5767 20964 7380 20992
rect 5767 20961 5779 20964
rect 5721 20955 5779 20961
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 8220 20992 8248 21032
rect 10594 21020 10600 21072
rect 10652 21060 10658 21072
rect 11790 21060 11796 21072
rect 10652 21032 11796 21060
rect 10652 21020 10658 21032
rect 11790 21020 11796 21032
rect 11848 21020 11854 21072
rect 8220 20964 8432 20992
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 8404 20924 8432 20964
rect 8478 20952 8484 21004
rect 8536 20952 8542 21004
rect 12176 20992 12204 21100
rect 13817 21097 13829 21100
rect 13863 21128 13875 21131
rect 16022 21128 16028 21140
rect 13863 21100 16028 21128
rect 13863 21097 13875 21100
rect 13817 21091 13875 21097
rect 16022 21088 16028 21100
rect 16080 21088 16086 21140
rect 16206 21088 16212 21140
rect 16264 21128 16270 21140
rect 24118 21128 24124 21140
rect 16264 21100 24124 21128
rect 16264 21088 16270 21100
rect 24118 21088 24124 21100
rect 24176 21088 24182 21140
rect 30650 21128 30656 21140
rect 25240 21100 30656 21128
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 14090 21060 14096 21072
rect 12308 21032 14096 21060
rect 12308 21020 12314 21032
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 16758 21060 16764 21072
rect 16316 21032 16764 21060
rect 9232 20964 9536 20992
rect 9232 20924 9260 20964
rect 7064 20896 8156 20924
rect 8404 20896 9260 20924
rect 7064 20884 7070 20896
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 2866 20856 2872 20868
rect 2823 20828 2872 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 8128 20856 8156 20896
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 9508 20924 9536 20964
rect 9646 20964 12204 20992
rect 9646 20924 9674 20964
rect 12526 20952 12532 21004
rect 12584 20952 12590 21004
rect 13725 20995 13783 21001
rect 13725 20961 13737 20995
rect 13771 20992 13783 20995
rect 13814 20992 13820 21004
rect 13771 20964 13820 20992
rect 13771 20961 13783 20964
rect 13725 20955 13783 20961
rect 13814 20952 13820 20964
rect 13872 20992 13878 21004
rect 14182 20992 14188 21004
rect 13872 20964 14188 20992
rect 13872 20952 13878 20964
rect 14182 20952 14188 20964
rect 14240 20992 14246 21004
rect 14458 20992 14464 21004
rect 14240 20964 14464 20992
rect 14240 20952 14246 20964
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 15102 20952 15108 21004
rect 15160 20952 15166 21004
rect 16316 20992 16344 21032
rect 16758 21020 16764 21032
rect 16816 21020 16822 21072
rect 21637 21063 21695 21069
rect 17604 21032 18920 21060
rect 17604 21001 17632 21032
rect 16132 20964 16344 20992
rect 16393 20995 16451 21001
rect 9508 20896 9674 20924
rect 10965 20927 11023 20933
rect 10965 20893 10977 20927
rect 11011 20924 11023 20927
rect 11146 20924 11152 20936
rect 11011 20896 11152 20924
rect 11011 20893 11023 20896
rect 10965 20887 11023 20893
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 12066 20884 12072 20936
rect 12124 20884 12130 20936
rect 15013 20927 15071 20933
rect 15013 20893 15025 20927
rect 15059 20924 15071 20927
rect 16132 20924 16160 20964
rect 16393 20961 16405 20995
rect 16439 20992 16451 20995
rect 17589 20995 17647 21001
rect 16439 20964 16804 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 15059 20896 16160 20924
rect 15059 20893 15071 20896
rect 15013 20887 15071 20893
rect 16206 20884 16212 20936
rect 16264 20884 16270 20936
rect 8205 20859 8263 20865
rect 8205 20856 8217 20859
rect 6946 20828 7420 20856
rect 8128 20828 8217 20856
rect 5169 20791 5227 20797
rect 5169 20757 5181 20791
rect 5215 20788 5227 20791
rect 6362 20788 6368 20800
rect 5215 20760 6368 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 6362 20748 6368 20760
rect 6420 20788 6426 20800
rect 7024 20788 7052 20828
rect 7392 20800 7420 20828
rect 8205 20825 8217 20828
rect 8251 20825 8263 20859
rect 8205 20819 8263 20825
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 10045 20859 10103 20865
rect 10045 20856 10057 20859
rect 8444 20828 10057 20856
rect 8444 20816 8450 20828
rect 10045 20825 10057 20828
rect 10091 20825 10103 20859
rect 10045 20819 10103 20825
rect 11330 20816 11336 20868
rect 11388 20816 11394 20868
rect 16482 20856 16488 20868
rect 14568 20828 16488 20856
rect 6420 20760 7052 20788
rect 6420 20748 6426 20760
rect 7190 20748 7196 20800
rect 7248 20748 7254 20800
rect 7374 20748 7380 20800
rect 7432 20788 7438 20800
rect 7469 20791 7527 20797
rect 7469 20788 7481 20791
rect 7432 20760 7481 20788
rect 7432 20748 7438 20760
rect 7469 20757 7481 20760
rect 7515 20757 7527 20791
rect 7469 20751 7527 20757
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 8110 20788 8116 20800
rect 7883 20760 8116 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 8297 20791 8355 20797
rect 8297 20757 8309 20791
rect 8343 20788 8355 20791
rect 10594 20788 10600 20800
rect 8343 20760 10600 20788
rect 8343 20757 8355 20760
rect 8297 20751 8355 20757
rect 10594 20748 10600 20760
rect 10652 20748 10658 20800
rect 11422 20748 11428 20800
rect 11480 20748 11486 20800
rect 14568 20797 14596 20828
rect 16482 20816 16488 20828
rect 16540 20816 16546 20868
rect 16776 20856 16804 20964
rect 17589 20961 17601 20995
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18601 20995 18659 21001
rect 18601 20992 18613 20995
rect 18012 20964 18613 20992
rect 18012 20952 18018 20964
rect 18601 20961 18613 20964
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 18782 20952 18788 21004
rect 18840 20952 18846 21004
rect 18892 20992 18920 21032
rect 21637 21029 21649 21063
rect 21683 21060 21695 21063
rect 21818 21060 21824 21072
rect 21683 21032 21824 21060
rect 21683 21029 21695 21032
rect 21637 21023 21695 21029
rect 21818 21020 21824 21032
rect 21876 21020 21882 21072
rect 24394 21060 24400 21072
rect 22066 21032 24400 21060
rect 19702 20992 19708 21004
rect 18892 20964 19708 20992
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 20254 20952 20260 21004
rect 20312 20992 20318 21004
rect 22066 20992 22094 21032
rect 24394 21020 24400 21032
rect 24452 21020 24458 21072
rect 20312 20964 22094 20992
rect 20312 20952 20318 20964
rect 22738 20952 22744 21004
rect 22796 20952 22802 21004
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20992 25191 20995
rect 25240 20992 25268 21100
rect 30650 21088 30656 21100
rect 30708 21088 30714 21140
rect 32493 21131 32551 21137
rect 32493 21097 32505 21131
rect 32539 21128 32551 21131
rect 32582 21128 32588 21140
rect 32539 21100 32588 21128
rect 32539 21097 32551 21100
rect 32493 21091 32551 21097
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 25958 21060 25964 21072
rect 25332 21032 25964 21060
rect 25332 21001 25360 21032
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 27614 21020 27620 21072
rect 27672 21060 27678 21072
rect 27672 21032 28580 21060
rect 27672 21020 27678 21032
rect 25179 20964 25268 20992
rect 25317 20995 25375 21001
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 25317 20961 25329 20995
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 25590 20952 25596 21004
rect 25648 20992 25654 21004
rect 26050 20992 26056 21004
rect 25648 20964 26056 20992
rect 25648 20952 25654 20964
rect 26050 20952 26056 20964
rect 26108 20992 26114 21004
rect 28350 20992 28356 21004
rect 26108 20964 28356 20992
rect 26108 20952 26114 20964
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 28552 21001 28580 21032
rect 28718 21020 28724 21072
rect 28776 21060 28782 21072
rect 36538 21060 36544 21072
rect 28776 21032 36544 21060
rect 28776 21020 28782 21032
rect 36538 21020 36544 21032
rect 36596 21020 36602 21072
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20961 28595 20995
rect 28537 20955 28595 20961
rect 30006 20952 30012 21004
rect 30064 20952 30070 21004
rect 17402 20884 17408 20936
rect 17460 20884 17466 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18874 20924 18880 20936
rect 18555 20896 18880 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 27614 20884 27620 20936
rect 27672 20924 27678 20936
rect 28261 20927 28319 20933
rect 27672 20896 27936 20924
rect 27672 20884 27678 20896
rect 16776 20828 19334 20856
rect 14553 20791 14611 20797
rect 14553 20757 14565 20791
rect 14599 20757 14611 20791
rect 14553 20751 14611 20757
rect 14921 20791 14979 20797
rect 14921 20757 14933 20791
rect 14967 20788 14979 20791
rect 15654 20788 15660 20800
rect 14967 20760 15660 20788
rect 14967 20757 14979 20760
rect 14921 20751 14979 20757
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 15746 20748 15752 20800
rect 15804 20748 15810 20800
rect 16117 20791 16175 20797
rect 16117 20757 16129 20791
rect 16163 20788 16175 20791
rect 16666 20788 16672 20800
rect 16163 20760 16672 20788
rect 16163 20757 16175 20760
rect 16117 20751 16175 20757
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17313 20791 17371 20797
rect 17313 20757 17325 20791
rect 17359 20788 17371 20791
rect 17770 20788 17776 20800
rect 17359 20760 17776 20788
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18322 20788 18328 20800
rect 18187 20760 18328 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18322 20748 18328 20760
rect 18380 20748 18386 20800
rect 19306 20788 19334 20828
rect 20714 20816 20720 20868
rect 20772 20816 20778 20868
rect 22465 20859 22523 20865
rect 22465 20825 22477 20859
rect 22511 20856 22523 20859
rect 23382 20856 23388 20868
rect 22511 20828 23388 20856
rect 22511 20825 22523 20828
rect 22465 20819 22523 20825
rect 23382 20816 23388 20828
rect 23440 20816 23446 20868
rect 23658 20816 23664 20868
rect 23716 20816 23722 20868
rect 25041 20859 25099 20865
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 26234 20856 26240 20868
rect 25087 20828 26240 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20825 26387 20859
rect 26329 20819 26387 20825
rect 20438 20788 20444 20800
rect 19306 20760 20444 20788
rect 20438 20748 20444 20760
rect 20496 20748 20502 20800
rect 20530 20748 20536 20800
rect 20588 20788 20594 20800
rect 21177 20791 21235 20797
rect 21177 20788 21189 20791
rect 20588 20760 21189 20788
rect 20588 20748 20594 20760
rect 21177 20757 21189 20760
rect 21223 20757 21235 20791
rect 21177 20751 21235 20757
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20788 22155 20791
rect 22186 20788 22192 20800
rect 22143 20760 22192 20788
rect 22143 20757 22155 20760
rect 22097 20751 22155 20757
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 22554 20748 22560 20800
rect 22612 20748 22618 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22704 20760 23305 20788
rect 22704 20748 22710 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 23293 20751 23351 20757
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 23753 20791 23811 20797
rect 23753 20788 23765 20791
rect 23532 20760 23765 20788
rect 23532 20748 23538 20760
rect 23753 20757 23765 20760
rect 23799 20757 23811 20791
rect 23753 20751 23811 20757
rect 24026 20748 24032 20800
rect 24084 20788 24090 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 24084 20760 24685 20788
rect 24084 20748 24090 20760
rect 24673 20757 24685 20760
rect 24719 20757 24731 20791
rect 24673 20751 24731 20757
rect 24762 20748 24768 20800
rect 24820 20788 24826 20800
rect 25777 20791 25835 20797
rect 25777 20788 25789 20791
rect 24820 20760 25789 20788
rect 24820 20748 24826 20760
rect 25777 20757 25789 20760
rect 25823 20788 25835 20791
rect 25866 20788 25872 20800
rect 25823 20760 25872 20788
rect 25823 20757 25835 20760
rect 25777 20751 25835 20757
rect 25866 20748 25872 20760
rect 25924 20748 25930 20800
rect 26344 20788 26372 20819
rect 26602 20816 26608 20868
rect 26660 20856 26666 20868
rect 27908 20856 27936 20896
rect 28261 20893 28273 20927
rect 28307 20924 28319 20927
rect 28442 20924 28448 20936
rect 28307 20896 28448 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28994 20884 29000 20936
rect 29052 20924 29058 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29052 20896 29745 20924
rect 29052 20884 29058 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 31849 20927 31907 20933
rect 31849 20924 31861 20927
rect 29733 20887 29791 20893
rect 29840 20896 31861 20924
rect 29840 20856 29868 20896
rect 31849 20893 31861 20896
rect 31895 20893 31907 20927
rect 31849 20887 31907 20893
rect 32677 20927 32735 20933
rect 32677 20893 32689 20927
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 30926 20856 30932 20868
rect 26660 20828 26818 20856
rect 27908 20828 29868 20856
rect 30300 20828 30932 20856
rect 26660 20816 26666 20828
rect 27614 20788 27620 20800
rect 26344 20760 27620 20788
rect 27614 20748 27620 20760
rect 27672 20748 27678 20800
rect 27801 20791 27859 20797
rect 27801 20757 27813 20791
rect 27847 20788 27859 20791
rect 27982 20788 27988 20800
rect 27847 20760 27988 20788
rect 27847 20757 27859 20760
rect 27801 20751 27859 20757
rect 27982 20748 27988 20760
rect 28040 20748 28046 20800
rect 28074 20748 28080 20800
rect 28132 20788 28138 20800
rect 28810 20788 28816 20800
rect 28132 20760 28816 20788
rect 28132 20748 28138 20760
rect 28810 20748 28816 20760
rect 28868 20788 28874 20800
rect 30300 20788 30328 20828
rect 30926 20816 30932 20828
rect 30984 20816 30990 20868
rect 31110 20816 31116 20868
rect 31168 20816 31174 20868
rect 31754 20816 31760 20868
rect 31812 20856 31818 20868
rect 32692 20856 32720 20887
rect 31812 20828 32720 20856
rect 31812 20816 31818 20828
rect 28868 20760 30328 20788
rect 28868 20748 28874 20760
rect 30374 20748 30380 20800
rect 30432 20788 30438 20800
rect 31205 20791 31263 20797
rect 31205 20788 31217 20791
rect 30432 20760 31217 20788
rect 30432 20748 30438 20760
rect 31205 20757 31217 20760
rect 31251 20757 31263 20791
rect 31205 20751 31263 20757
rect 31938 20748 31944 20800
rect 31996 20748 32002 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 11422 20584 11428 20596
rect 4396 20556 11428 20584
rect 4396 20544 4402 20556
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13035 20556 15792 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 3878 20476 3884 20528
rect 3936 20516 3942 20528
rect 8757 20519 8815 20525
rect 3936 20488 7052 20516
rect 3936 20476 3942 20488
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 4062 20448 4068 20460
rect 3651 20420 4068 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 4062 20408 4068 20420
rect 4120 20408 4126 20460
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20448 5687 20451
rect 5675 20420 6040 20448
rect 5675 20417 5687 20420
rect 5629 20411 5687 20417
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5721 20383 5779 20389
rect 5721 20349 5733 20383
rect 5767 20349 5779 20383
rect 5721 20343 5779 20349
rect 5736 20312 5764 20343
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 6012 20380 6040 20420
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6144 20420 6561 20448
rect 6144 20408 6150 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6822 20380 6828 20392
rect 6012 20352 6828 20380
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7024 20389 7052 20488
rect 8757 20485 8769 20519
rect 8803 20516 8815 20519
rect 9950 20516 9956 20528
rect 8803 20488 9956 20516
rect 8803 20485 8815 20488
rect 8757 20479 8815 20485
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 11146 20516 11152 20528
rect 10902 20488 11152 20516
rect 11146 20476 11152 20488
rect 11204 20476 11210 20528
rect 12526 20476 12532 20528
rect 12584 20516 12590 20528
rect 13538 20516 13544 20528
rect 12584 20488 13544 20516
rect 12584 20476 12590 20488
rect 13538 20476 13544 20488
rect 13596 20516 13602 20528
rect 13596 20488 13768 20516
rect 13596 20476 13602 20488
rect 7374 20408 7380 20460
rect 7432 20448 7438 20460
rect 8389 20451 8447 20457
rect 8389 20448 8401 20451
rect 7432 20420 8401 20448
rect 7432 20408 7438 20420
rect 8389 20417 8401 20420
rect 8435 20448 8447 20451
rect 8938 20448 8944 20460
rect 8435 20420 8944 20448
rect 8435 20417 8447 20420
rect 8389 20411 8447 20417
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 12802 20448 12808 20460
rect 11848 20420 12808 20448
rect 11848 20408 11854 20420
rect 12802 20408 12808 20420
rect 12860 20408 12866 20460
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 13630 20448 13636 20460
rect 13495 20420 13636 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 9398 20340 9404 20392
rect 9456 20340 9462 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 9732 20352 11100 20380
rect 9732 20340 9738 20352
rect 6086 20312 6092 20324
rect 5736 20284 6092 20312
rect 6086 20272 6092 20284
rect 6144 20272 6150 20324
rect 7374 20272 7380 20324
rect 7432 20312 7438 20324
rect 8941 20315 8999 20321
rect 8941 20312 8953 20315
rect 7432 20284 8953 20312
rect 7432 20272 7438 20284
rect 8941 20281 8953 20284
rect 8987 20281 8999 20315
rect 11072 20312 11100 20352
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 12250 20380 12256 20392
rect 11204 20352 12256 20380
rect 11204 20340 11210 20352
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12526 20380 12532 20392
rect 12483 20352 12532 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12526 20340 12532 20352
rect 12584 20380 12590 20392
rect 12912 20380 12940 20411
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 13740 20457 13768 20488
rect 14458 20476 14464 20528
rect 14516 20476 14522 20528
rect 15764 20516 15792 20556
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17000 20556 17509 20584
rect 17000 20544 17006 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 17497 20547 17555 20553
rect 18509 20587 18567 20593
rect 18509 20553 18521 20587
rect 18555 20553 18567 20587
rect 18509 20547 18567 20553
rect 18524 20516 18552 20547
rect 18874 20544 18880 20596
rect 18932 20544 18938 20596
rect 18969 20587 19027 20593
rect 18969 20553 18981 20587
rect 19015 20584 19027 20587
rect 19058 20584 19064 20596
rect 19015 20556 19064 20584
rect 19015 20553 19027 20556
rect 18969 20547 19027 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19484 20556 22784 20584
rect 19484 20544 19490 20556
rect 15764 20488 18552 20516
rect 18800 20488 19012 20516
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 16022 20408 16028 20460
rect 16080 20408 16086 20460
rect 17405 20451 17463 20457
rect 17405 20448 17417 20451
rect 16132 20420 17417 20448
rect 12584 20352 12940 20380
rect 13173 20383 13231 20389
rect 12584 20340 12590 20352
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13219 20352 13860 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13446 20312 13452 20324
rect 11072 20284 13452 20312
rect 8941 20275 8999 20281
rect 13446 20272 13452 20284
rect 13504 20272 13510 20324
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 7098 20244 7104 20256
rect 5307 20216 7104 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 9030 20204 9036 20256
rect 9088 20244 9094 20256
rect 10134 20244 10140 20256
rect 9088 20216 10140 20244
rect 9088 20204 9094 20216
rect 10134 20204 10140 20216
rect 10192 20244 10198 20256
rect 10870 20244 10876 20256
rect 10192 20216 10876 20244
rect 10192 20204 10198 20216
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 11882 20204 11888 20256
rect 11940 20204 11946 20256
rect 12529 20247 12587 20253
rect 12529 20213 12541 20247
rect 12575 20244 12587 20247
rect 12710 20244 12716 20256
rect 12575 20216 12716 20244
rect 12575 20213 12587 20216
rect 12529 20207 12587 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13630 20204 13636 20256
rect 13688 20204 13694 20256
rect 13832 20244 13860 20352
rect 13998 20340 14004 20392
rect 14056 20340 14062 20392
rect 14642 20340 14648 20392
rect 14700 20380 14706 20392
rect 16132 20380 16160 20420
rect 17405 20417 17417 20420
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 17494 20408 17500 20460
rect 17552 20448 17558 20460
rect 18800 20448 18828 20488
rect 17552 20420 18828 20448
rect 18984 20448 19012 20488
rect 18984 20420 19104 20448
rect 17552 20408 17558 20420
rect 14700 20352 16160 20380
rect 16761 20383 16819 20389
rect 14700 20340 14706 20352
rect 16761 20349 16773 20383
rect 16807 20380 16819 20383
rect 17589 20383 17647 20389
rect 16807 20352 17540 20380
rect 16807 20349 16819 20352
rect 16761 20343 16819 20349
rect 17126 20312 17132 20324
rect 15028 20284 17132 20312
rect 15028 20244 15056 20284
rect 17126 20272 17132 20284
rect 17184 20272 17190 20324
rect 13832 20216 15056 20244
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 17037 20247 17095 20253
rect 17037 20244 17049 20247
rect 16816 20216 17049 20244
rect 16816 20204 16822 20216
rect 17037 20213 17049 20216
rect 17083 20213 17095 20247
rect 17512 20244 17540 20352
rect 17589 20349 17601 20383
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 17604 20312 17632 20343
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18874 20380 18880 20392
rect 18012 20352 18880 20380
rect 18012 20340 18018 20352
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 19076 20389 19104 20420
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19610 20448 19616 20460
rect 19484 20420 19616 20448
rect 19484 20408 19490 20420
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 19720 20457 19748 20556
rect 20714 20476 20720 20528
rect 20772 20476 20778 20528
rect 22002 20476 22008 20528
rect 22060 20476 22066 20528
rect 22756 20525 22784 20556
rect 23382 20544 23388 20596
rect 23440 20544 23446 20596
rect 23658 20544 23664 20596
rect 23716 20584 23722 20596
rect 24762 20584 24768 20596
rect 23716 20556 24768 20584
rect 23716 20544 23722 20556
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 27246 20544 27252 20596
rect 27304 20584 27310 20596
rect 27525 20587 27583 20593
rect 27525 20584 27537 20587
rect 27304 20556 27537 20584
rect 27304 20544 27310 20556
rect 27525 20553 27537 20556
rect 27571 20553 27583 20587
rect 27525 20547 27583 20553
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 28534 20584 28540 20596
rect 27663 20556 28540 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 22741 20519 22799 20525
rect 22741 20485 22753 20519
rect 22787 20485 22799 20519
rect 22741 20479 22799 20485
rect 25866 20476 25872 20528
rect 25924 20516 25930 20528
rect 27264 20516 27292 20544
rect 25924 20488 27292 20516
rect 27540 20516 27568 20547
rect 28534 20544 28540 20556
rect 28592 20544 28598 20596
rect 31021 20587 31079 20593
rect 31021 20553 31033 20587
rect 31067 20584 31079 20587
rect 34974 20584 34980 20596
rect 31067 20556 34980 20584
rect 31067 20553 31079 20556
rect 31021 20547 31079 20553
rect 34974 20544 34980 20556
rect 35032 20544 35038 20596
rect 27798 20516 27804 20528
rect 27540 20488 27804 20516
rect 25924 20476 25930 20488
rect 27798 20476 27804 20488
rect 27856 20476 27862 20528
rect 28629 20519 28687 20525
rect 28629 20485 28641 20519
rect 28675 20516 28687 20519
rect 28902 20516 28908 20528
rect 28675 20488 28908 20516
rect 28675 20485 28687 20488
rect 28629 20479 28687 20485
rect 28902 20476 28908 20488
rect 28960 20476 28966 20528
rect 29086 20476 29092 20528
rect 29144 20476 29150 20528
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 23348 20420 24317 20448
rect 23348 20408 23354 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 26421 20451 26479 20457
rect 26421 20448 26433 20451
rect 25714 20434 26433 20448
rect 24305 20411 24363 20417
rect 25700 20420 26433 20434
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20380 19119 20383
rect 19981 20383 20039 20389
rect 19107 20352 19748 20380
rect 19107 20349 19119 20352
rect 19061 20343 19119 20349
rect 19610 20312 19616 20324
rect 17604 20284 19616 20312
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 17954 20244 17960 20256
rect 17512 20216 17960 20244
rect 17037 20207 17095 20213
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 18233 20247 18291 20253
rect 18233 20213 18245 20247
rect 18279 20244 18291 20247
rect 18690 20244 18696 20256
rect 18279 20216 18696 20244
rect 18279 20213 18291 20216
rect 18233 20207 18291 20213
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 19242 20244 19248 20256
rect 18932 20216 19248 20244
rect 18932 20204 18938 20216
rect 19242 20204 19248 20216
rect 19300 20204 19306 20256
rect 19720 20244 19748 20352
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20622 20380 20628 20392
rect 20027 20352 20628 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 24026 20340 24032 20392
rect 24084 20340 24090 20392
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 24670 20380 24676 20392
rect 24627 20352 24676 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 24670 20340 24676 20352
rect 24728 20340 24734 20392
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25700 20380 25728 20420
rect 26421 20417 26433 20420
rect 26467 20448 26479 20451
rect 26510 20448 26516 20460
rect 26467 20420 26516 20448
rect 26467 20417 26479 20420
rect 26421 20411 26479 20417
rect 26510 20408 26516 20420
rect 26568 20448 26574 20460
rect 26697 20451 26755 20457
rect 26697 20448 26709 20451
rect 26568 20420 26709 20448
rect 26568 20408 26574 20420
rect 26697 20417 26709 20420
rect 26743 20417 26755 20451
rect 26697 20411 26755 20417
rect 28350 20408 28356 20460
rect 28408 20408 28414 20460
rect 30929 20451 30987 20457
rect 30929 20448 30941 20451
rect 29840 20420 30941 20448
rect 25188 20352 25728 20380
rect 25188 20340 25194 20352
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 26016 20352 26065 20380
rect 26016 20340 26022 20352
rect 26053 20349 26065 20352
rect 26099 20380 26111 20383
rect 27709 20383 27767 20389
rect 27709 20380 27721 20383
rect 26099 20352 27721 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 27709 20349 27721 20352
rect 27755 20349 27767 20383
rect 29840 20380 29868 20420
rect 30929 20417 30941 20420
rect 30975 20448 30987 20451
rect 31573 20451 31631 20457
rect 31573 20448 31585 20451
rect 30975 20420 31585 20448
rect 30975 20417 30987 20420
rect 30929 20411 30987 20417
rect 31573 20417 31585 20420
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 27709 20343 27767 20349
rect 28460 20352 29868 20380
rect 26326 20272 26332 20324
rect 26384 20312 26390 20324
rect 26384 20284 27384 20312
rect 26384 20272 26390 20284
rect 21453 20247 21511 20253
rect 21453 20244 21465 20247
rect 19720 20216 21465 20244
rect 21453 20213 21465 20216
rect 21499 20213 21511 20247
rect 21453 20207 21511 20213
rect 22554 20204 22560 20256
rect 22612 20244 22618 20256
rect 27157 20247 27215 20253
rect 27157 20244 27169 20247
rect 22612 20216 27169 20244
rect 22612 20204 22618 20216
rect 27157 20213 27169 20216
rect 27203 20213 27215 20247
rect 27356 20244 27384 20284
rect 27430 20272 27436 20324
rect 27488 20312 27494 20324
rect 28460 20312 28488 20352
rect 30006 20340 30012 20392
rect 30064 20380 30070 20392
rect 31113 20383 31171 20389
rect 31113 20380 31125 20383
rect 30064 20352 31125 20380
rect 30064 20340 30070 20352
rect 31113 20349 31125 20352
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 27488 20284 28488 20312
rect 27488 20272 27494 20284
rect 30101 20247 30159 20253
rect 30101 20244 30113 20247
rect 27356 20216 30113 20244
rect 27157 20207 27215 20213
rect 30101 20213 30113 20216
rect 30147 20213 30159 20247
rect 30101 20207 30159 20213
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 30561 20247 30619 20253
rect 30561 20244 30573 20247
rect 30248 20216 30573 20244
rect 30248 20204 30254 20216
rect 30561 20213 30573 20216
rect 30607 20213 30619 20247
rect 30561 20207 30619 20213
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 4338 20040 4344 20052
rect 1780 20012 4344 20040
rect 1780 19845 1808 20012
rect 4338 20000 4344 20012
rect 4396 20000 4402 20052
rect 5442 20040 5448 20052
rect 4540 20012 5448 20040
rect 4540 19913 4568 20012
rect 5442 20000 5448 20012
rect 5500 20040 5506 20052
rect 8294 20040 8300 20052
rect 5500 20012 8300 20040
rect 5500 20000 5506 20012
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19873 4583 19907
rect 4525 19867 4583 19873
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19904 4859 19907
rect 6362 19904 6368 19916
rect 4847 19876 6368 19904
rect 4847 19873 4859 19876
rect 4801 19867 4859 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 6748 19913 6776 20012
rect 8294 20000 8300 20012
rect 8352 20040 8358 20052
rect 9398 20040 9404 20052
rect 8352 20012 9404 20040
rect 8352 20000 8358 20012
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 10870 20000 10876 20052
rect 10928 20000 10934 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11149 20043 11207 20049
rect 11149 20040 11161 20043
rect 11112 20012 11161 20040
rect 11112 20000 11118 20012
rect 11149 20009 11161 20012
rect 11195 20009 11207 20043
rect 11149 20003 11207 20009
rect 11517 20043 11575 20049
rect 11517 20009 11529 20043
rect 11563 20040 11575 20043
rect 11790 20040 11796 20052
rect 11563 20012 11796 20040
rect 11563 20009 11575 20012
rect 11517 20003 11575 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12989 20043 13047 20049
rect 12989 20009 13001 20043
rect 13035 20040 13047 20043
rect 13354 20040 13360 20052
rect 13035 20012 13360 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 13998 20000 14004 20052
rect 14056 20040 14062 20052
rect 15010 20040 15016 20052
rect 14056 20012 15016 20040
rect 14056 20000 14062 20012
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19886 20040 19892 20052
rect 18739 20012 19892 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19886 20000 19892 20012
rect 19944 20000 19950 20052
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 23382 20040 23388 20052
rect 21232 20012 23388 20040
rect 21232 20000 21238 20012
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 30745 20043 30803 20049
rect 30745 20040 30757 20043
rect 25148 20012 30757 20040
rect 12434 19972 12440 19984
rect 10704 19944 12440 19972
rect 6733 19907 6791 19913
rect 6733 19873 6745 19907
rect 6779 19873 6791 19907
rect 6733 19867 6791 19873
rect 7009 19907 7067 19913
rect 7009 19873 7021 19907
rect 7055 19904 7067 19907
rect 9030 19904 9036 19916
rect 7055 19876 9036 19904
rect 7055 19873 7067 19876
rect 7009 19867 7067 19873
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 10704 19904 10732 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 12802 19932 12808 19984
rect 12860 19972 12866 19984
rect 14366 19972 14372 19984
rect 12860 19944 14372 19972
rect 12860 19932 12866 19944
rect 14366 19932 14372 19944
rect 14424 19932 14430 19984
rect 16945 19975 17003 19981
rect 16945 19941 16957 19975
rect 16991 19972 17003 19975
rect 17770 19972 17776 19984
rect 16991 19944 17776 19972
rect 16991 19941 17003 19944
rect 16945 19935 17003 19941
rect 17770 19932 17776 19944
rect 17828 19932 17834 19984
rect 20254 19972 20260 19984
rect 19536 19944 20260 19972
rect 9171 19876 10732 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 12342 19864 12348 19916
rect 12400 19864 12406 19916
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13679 19876 14841 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14829 19873 14841 19876
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 18966 19904 18972 19916
rect 17911 19876 18972 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 18966 19864 18972 19876
rect 19024 19904 19030 19916
rect 19242 19904 19248 19916
rect 19024 19876 19248 19904
rect 19024 19864 19030 19876
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19805 1823 19839
rect 1765 19799 1823 19805
rect 10502 19796 10508 19848
rect 10560 19836 10566 19848
rect 11054 19836 11060 19848
rect 10560 19808 11060 19836
rect 10560 19796 10566 19808
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 12158 19796 12164 19848
rect 12216 19796 12222 19848
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 14458 19836 14464 19848
rect 12299 19808 14464 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 18322 19836 18328 19848
rect 17727 19808 18328 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19058 19836 19064 19848
rect 18923 19808 19064 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 2777 19771 2835 19777
rect 2777 19737 2789 19771
rect 2823 19768 2835 19771
rect 2866 19768 2872 19780
rect 2823 19740 2872 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 6178 19768 6184 19780
rect 6026 19740 6184 19768
rect 6178 19728 6184 19740
rect 6236 19768 6242 19780
rect 7466 19768 7472 19780
rect 6236 19740 7472 19768
rect 6236 19728 6242 19740
rect 7466 19728 7472 19740
rect 7524 19728 7530 19780
rect 9401 19771 9459 19777
rect 9401 19737 9413 19771
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 3694 19660 3700 19712
rect 3752 19700 3758 19712
rect 4246 19700 4252 19712
rect 3752 19672 4252 19700
rect 3752 19660 3758 19672
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 6273 19703 6331 19709
rect 6273 19669 6285 19703
rect 6319 19700 6331 19703
rect 7834 19700 7840 19712
rect 6319 19672 7840 19700
rect 6319 19669 6331 19672
rect 6273 19663 6331 19669
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 8481 19703 8539 19709
rect 8481 19700 8493 19703
rect 8352 19672 8493 19700
rect 8352 19660 8358 19672
rect 8481 19669 8493 19672
rect 8527 19669 8539 19703
rect 9416 19700 9444 19731
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 12618 19768 12624 19780
rect 11020 19740 12624 19768
rect 11020 19728 11026 19740
rect 12618 19728 12624 19740
rect 12676 19728 12682 19780
rect 12802 19728 12808 19780
rect 12860 19768 12866 19780
rect 13357 19771 13415 19777
rect 13357 19768 13369 19771
rect 12860 19740 13369 19768
rect 12860 19728 12866 19740
rect 13357 19737 13369 19740
rect 13403 19737 13415 19771
rect 13357 19731 13415 19737
rect 13449 19771 13507 19777
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 13495 19740 15240 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 11146 19700 11152 19712
rect 9416 19672 11152 19700
rect 8481 19663 8539 19669
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11790 19660 11796 19712
rect 11848 19660 11854 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 13630 19700 13636 19712
rect 12768 19672 13636 19700
rect 12768 19660 12774 19672
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 13906 19660 13912 19712
rect 13964 19660 13970 19712
rect 14182 19660 14188 19712
rect 14240 19660 14246 19712
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14461 19703 14519 19709
rect 14461 19700 14473 19703
rect 14424 19672 14473 19700
rect 14424 19660 14430 19672
rect 14461 19669 14473 19672
rect 14507 19700 14519 19703
rect 14826 19700 14832 19712
rect 14507 19672 14832 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 15212 19700 15240 19740
rect 15286 19728 15292 19780
rect 15344 19728 15350 19780
rect 16224 19740 18368 19768
rect 16224 19700 16252 19740
rect 18340 19712 18368 19740
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 19536 19768 19564 19944
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 22922 19932 22928 19984
rect 22980 19972 22986 19984
rect 24673 19975 24731 19981
rect 24673 19972 24685 19975
rect 22980 19944 24685 19972
rect 22980 19932 22986 19944
rect 24673 19941 24685 19944
rect 24719 19941 24731 19975
rect 24673 19935 24731 19941
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 20530 19904 20536 19916
rect 19668 19876 20536 19904
rect 19668 19864 19674 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 23842 19904 23848 19916
rect 22020 19876 23848 19904
rect 19702 19796 19708 19848
rect 19760 19836 19766 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 19760 19808 20269 19836
rect 19760 19796 19766 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 19024 19740 19564 19768
rect 19613 19771 19671 19777
rect 19024 19728 19030 19740
rect 19613 19737 19625 19771
rect 19659 19768 19671 19771
rect 19978 19768 19984 19780
rect 19659 19740 19984 19768
rect 19659 19737 19671 19740
rect 19613 19731 19671 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 20732 19740 21022 19768
rect 20732 19712 20760 19740
rect 15212 19672 16252 19700
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 16390 19700 16396 19712
rect 16347 19672 16396 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 16761 19703 16819 19709
rect 16761 19669 16773 19703
rect 16807 19700 16819 19703
rect 16942 19700 16948 19712
rect 16807 19672 16948 19700
rect 16807 19669 16819 19672
rect 16761 19663 16819 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 17586 19660 17592 19712
rect 17644 19660 17650 19712
rect 18322 19660 18328 19712
rect 18380 19660 18386 19712
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19886 19700 19892 19712
rect 19751 19672 19892 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 20714 19660 20720 19712
rect 20772 19660 20778 19712
rect 21450 19660 21456 19712
rect 21508 19700 21514 19712
rect 22020 19709 22048 19876
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 25148 19913 25176 20012
rect 30745 20009 30757 20012
rect 30791 20009 30803 20043
rect 48314 20040 48320 20052
rect 30745 20003 30803 20009
rect 30852 20012 48320 20040
rect 27614 19932 27620 19984
rect 27672 19932 27678 19984
rect 29730 19932 29736 19984
rect 29788 19932 29794 19984
rect 30466 19932 30472 19984
rect 30524 19932 30530 19984
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 25317 19907 25375 19913
rect 25317 19873 25329 19907
rect 25363 19904 25375 19907
rect 26142 19904 26148 19916
rect 25363 19876 26148 19904
rect 25363 19873 25375 19876
rect 25317 19867 25375 19873
rect 26142 19864 26148 19876
rect 26200 19864 26206 19916
rect 27706 19864 27712 19916
rect 27764 19904 27770 19916
rect 28353 19907 28411 19913
rect 28353 19904 28365 19907
rect 27764 19876 28365 19904
rect 27764 19864 27770 19876
rect 28353 19873 28365 19876
rect 28399 19873 28411 19907
rect 28353 19867 28411 19873
rect 28626 19864 28632 19916
rect 28684 19864 28690 19916
rect 30852 19904 30880 20012
rect 48314 20000 48320 20012
rect 48372 20000 48378 20052
rect 28966 19876 30880 19904
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19836 22615 19839
rect 25498 19836 25504 19848
rect 22603 19808 25504 19836
rect 22603 19805 22615 19808
rect 22557 19799 22615 19805
rect 25498 19796 25504 19808
rect 25556 19796 25562 19848
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 28966 19836 28994 19876
rect 31294 19864 31300 19916
rect 31352 19864 31358 19916
rect 27580 19808 28994 19836
rect 27580 19796 27586 19808
rect 29914 19796 29920 19848
rect 29972 19796 29978 19848
rect 30466 19836 30472 19848
rect 30024 19808 30472 19836
rect 23753 19771 23811 19777
rect 23753 19737 23765 19771
rect 23799 19768 23811 19771
rect 24026 19768 24032 19780
rect 23799 19740 24032 19768
rect 23799 19737 23811 19740
rect 23753 19731 23811 19737
rect 24026 19728 24032 19740
rect 24084 19768 24090 19780
rect 25222 19768 25228 19780
rect 24084 19740 25228 19768
rect 24084 19728 24090 19740
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 25682 19728 25688 19780
rect 25740 19768 25746 19780
rect 26145 19771 26203 19777
rect 26145 19768 26157 19771
rect 25740 19740 26157 19768
rect 25740 19728 25746 19740
rect 26145 19737 26157 19740
rect 26191 19737 26203 19771
rect 26145 19731 26203 19737
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 28350 19728 28356 19780
rect 28408 19768 28414 19780
rect 30024 19768 30052 19808
rect 30466 19796 30472 19808
rect 30524 19836 30530 19848
rect 31113 19839 31171 19845
rect 31113 19836 31125 19839
rect 30524 19808 31125 19836
rect 30524 19796 30530 19808
rect 31113 19805 31125 19808
rect 31159 19805 31171 19839
rect 31113 19799 31171 19805
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19836 31263 19839
rect 34606 19836 34612 19848
rect 31251 19808 34612 19836
rect 31251 19805 31263 19808
rect 31205 19799 31263 19805
rect 34606 19796 34612 19808
rect 34664 19796 34670 19848
rect 28408 19740 30052 19768
rect 28408 19728 28414 19740
rect 22005 19703 22063 19709
rect 22005 19700 22017 19703
rect 21508 19672 22017 19700
rect 21508 19660 21514 19672
rect 22005 19669 22017 19672
rect 22051 19669 22063 19703
rect 22005 19663 22063 19669
rect 22278 19660 22284 19712
rect 22336 19700 22342 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 22336 19672 22661 19700
rect 22336 19660 22342 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 22649 19663 22707 19669
rect 23290 19660 23296 19712
rect 23348 19660 23354 19712
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 25038 19660 25044 19712
rect 25096 19660 25102 19712
rect 27706 19660 27712 19712
rect 27764 19700 27770 19712
rect 27893 19703 27951 19709
rect 27893 19700 27905 19703
rect 27764 19672 27905 19700
rect 27764 19660 27770 19672
rect 27893 19669 27905 19672
rect 27939 19700 27951 19703
rect 29086 19700 29092 19712
rect 27939 19672 29092 19700
rect 27939 19669 27951 19672
rect 27893 19663 27951 19669
rect 29086 19660 29092 19672
rect 29144 19660 29150 19712
rect 30282 19660 30288 19712
rect 30340 19660 30346 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 4890 19496 4896 19508
rect 2746 19468 4896 19496
rect 2746 19428 2774 19468
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 5261 19499 5319 19505
rect 5261 19465 5273 19499
rect 5307 19465 5319 19499
rect 5261 19459 5319 19465
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 6454 19496 6460 19508
rect 5767 19468 6460 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 1780 19400 2774 19428
rect 1780 19369 1808 19400
rect 3510 19388 3516 19440
rect 3568 19428 3574 19440
rect 4341 19431 4399 19437
rect 4341 19428 4353 19431
rect 3568 19400 4353 19428
rect 3568 19388 3574 19400
rect 4341 19397 4353 19400
rect 4387 19397 4399 19431
rect 4341 19391 4399 19397
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 3694 19360 3700 19372
rect 3651 19332 3700 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 3694 19320 3700 19332
rect 3752 19320 3758 19372
rect 4522 19320 4528 19372
rect 4580 19360 4586 19372
rect 4890 19360 4896 19372
rect 4580 19332 4896 19360
rect 4580 19320 4586 19332
rect 4890 19320 4896 19332
rect 4948 19320 4954 19372
rect 5276 19360 5304 19459
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 10318 19496 10324 19508
rect 6840 19468 10324 19496
rect 5629 19431 5687 19437
rect 5629 19397 5641 19431
rect 5675 19428 5687 19431
rect 6840 19428 6868 19468
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 10410 19456 10416 19508
rect 10468 19456 10474 19508
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 10962 19496 10968 19508
rect 10919 19468 10968 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 14550 19496 14556 19508
rect 11992 19468 14556 19496
rect 11992 19440 12020 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 18325 19499 18383 19505
rect 14884 19468 18000 19496
rect 14884 19456 14890 19468
rect 5675 19400 6868 19428
rect 5675 19397 5687 19400
rect 5629 19391 5687 19397
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 7469 19431 7527 19437
rect 7469 19428 7481 19431
rect 6972 19400 7481 19428
rect 6972 19388 6978 19400
rect 7469 19397 7481 19400
rect 7515 19397 7527 19431
rect 7469 19391 7527 19397
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 7616 19400 9321 19428
rect 7616 19388 7622 19400
rect 9309 19397 9321 19400
rect 9355 19397 9367 19431
rect 9309 19391 9367 19397
rect 9950 19388 9956 19440
rect 10008 19428 10014 19440
rect 10137 19431 10195 19437
rect 10137 19428 10149 19431
rect 10008 19400 10149 19428
rect 10008 19388 10014 19400
rect 10137 19397 10149 19400
rect 10183 19428 10195 19431
rect 10686 19428 10692 19440
rect 10183 19400 10692 19428
rect 10183 19397 10195 19400
rect 10137 19391 10195 19397
rect 10686 19388 10692 19400
rect 10744 19388 10750 19440
rect 11974 19428 11980 19440
rect 11716 19400 11980 19428
rect 6454 19360 6460 19372
rect 5276 19332 6460 19360
rect 6454 19320 6460 19332
rect 6512 19320 6518 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 8662 19360 8668 19372
rect 8619 19332 8668 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 11716 19369 11744 19400
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 14182 19428 14188 19440
rect 13202 19400 14188 19428
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 14277 19431 14335 19437
rect 14277 19397 14289 19431
rect 14323 19428 14335 19431
rect 14366 19428 14372 19440
rect 14323 19400 14372 19428
rect 14323 19397 14335 19400
rect 14277 19391 14335 19397
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 10367 19332 10793 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10781 19329 10793 19332
rect 10827 19360 10839 19363
rect 11701 19363 11759 19369
rect 10827 19332 11100 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 11072 19304 11100 19332
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19292 5963 19295
rect 7190 19292 7196 19304
rect 5951 19264 7196 19292
rect 5951 19261 5963 19264
rect 5905 19255 5963 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 9732 19264 10977 19292
rect 9732 19252 9738 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 11054 19252 11060 19304
rect 11112 19252 11118 19304
rect 11977 19295 12035 19301
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 12023 19264 13032 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 4522 19184 4528 19236
rect 4580 19224 4586 19236
rect 13004 19224 13032 19264
rect 13446 19252 13452 19304
rect 13504 19252 13510 19304
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 14292 19292 14320 19391
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 14458 19388 14464 19440
rect 14516 19428 14522 19440
rect 17972 19428 18000 19468
rect 18325 19465 18337 19499
rect 18371 19496 18383 19499
rect 18506 19496 18512 19508
rect 18371 19468 18512 19496
rect 18371 19465 18383 19468
rect 18325 19459 18383 19465
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 19300 19468 21465 19496
rect 19300 19456 19306 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 23290 19496 23296 19508
rect 22419 19468 23296 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 23566 19456 23572 19508
rect 23624 19496 23630 19508
rect 23661 19499 23719 19505
rect 23661 19496 23673 19499
rect 23624 19468 23673 19496
rect 23624 19456 23630 19468
rect 23661 19465 23673 19468
rect 23707 19465 23719 19499
rect 23661 19459 23719 19465
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26421 19499 26479 19505
rect 26421 19496 26433 19499
rect 26292 19468 26433 19496
rect 26292 19456 26298 19468
rect 26421 19465 26433 19468
rect 26467 19465 26479 19499
rect 26421 19459 26479 19465
rect 26602 19456 26608 19508
rect 26660 19496 26666 19508
rect 30374 19496 30380 19508
rect 26660 19468 30380 19496
rect 26660 19456 26666 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 30469 19499 30527 19505
rect 30469 19465 30481 19499
rect 30515 19496 30527 19499
rect 30515 19468 31754 19496
rect 30515 19465 30527 19468
rect 30469 19459 30527 19465
rect 20070 19428 20076 19440
rect 14516 19400 17908 19428
rect 17972 19400 20076 19428
rect 14516 19388 14522 19400
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14476 19332 14749 19360
rect 14476 19304 14504 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 15838 19360 15844 19372
rect 15703 19332 15844 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 15838 19320 15844 19332
rect 15896 19360 15902 19372
rect 16022 19360 16028 19372
rect 15896 19332 16028 19360
rect 15896 19320 15902 19332
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 16485 19363 16543 19369
rect 16485 19360 16497 19363
rect 16224 19332 16497 19360
rect 16224 19304 16252 19332
rect 16485 19329 16497 19332
rect 16531 19360 16543 19363
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16531 19332 16773 19360
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 16761 19329 16773 19332
rect 16807 19360 16819 19363
rect 17405 19363 17463 19369
rect 16807 19332 16988 19360
rect 16807 19329 16819 19332
rect 16761 19323 16819 19329
rect 13964 19264 14320 19292
rect 13964 19252 13970 19264
rect 14458 19252 14464 19304
rect 14516 19252 14522 19304
rect 14826 19252 14832 19304
rect 14884 19292 14890 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14884 19264 14933 19292
rect 14884 19252 14890 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15010 19252 15016 19304
rect 15068 19292 15074 19304
rect 15068 19264 15976 19292
rect 15068 19252 15074 19264
rect 13262 19224 13268 19236
rect 4580 19196 10272 19224
rect 13004 19196 13268 19224
rect 4580 19184 4586 19196
rect 5442 19116 5448 19168
rect 5500 19156 5506 19168
rect 6546 19156 6552 19168
rect 5500 19128 6552 19156
rect 5500 19116 5506 19128
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 10244 19156 10272 19196
rect 13262 19184 13268 19196
rect 13320 19184 13326 19236
rect 13372 19196 14320 19224
rect 13372 19156 13400 19196
rect 10244 19128 13400 19156
rect 13725 19159 13783 19165
rect 13725 19125 13737 19159
rect 13771 19156 13783 19159
rect 13906 19156 13912 19168
rect 13771 19128 13912 19156
rect 13771 19125 13783 19128
rect 13725 19119 13783 19125
rect 13906 19116 13912 19128
rect 13964 19156 13970 19168
rect 14001 19159 14059 19165
rect 14001 19156 14013 19159
rect 13964 19128 14013 19156
rect 13964 19116 13970 19128
rect 14001 19125 14013 19128
rect 14047 19125 14059 19159
rect 14292 19156 14320 19196
rect 14366 19184 14372 19236
rect 14424 19184 14430 19236
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 14476 19196 15853 19224
rect 14476 19156 14504 19196
rect 15841 19193 15853 19196
rect 15887 19193 15899 19227
rect 15948 19224 15976 19264
rect 16206 19252 16212 19304
rect 16264 19252 16270 19304
rect 16960 19301 16988 19332
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 17770 19360 17776 19372
rect 17451 19332 17776 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19292 17003 19295
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 16991 19264 17141 19292
rect 16991 19261 17003 19264
rect 16945 19255 17003 19261
rect 17129 19261 17141 19264
rect 17175 19292 17187 19295
rect 17678 19292 17684 19304
rect 17175 19264 17684 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17678 19252 17684 19264
rect 17736 19252 17742 19304
rect 17880 19292 17908 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20714 19388 20720 19440
rect 20772 19388 20778 19440
rect 22465 19431 22523 19437
rect 22465 19397 22477 19431
rect 22511 19428 22523 19431
rect 22646 19428 22652 19440
rect 22511 19400 22652 19428
rect 22511 19397 22523 19400
rect 22465 19391 22523 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 23109 19431 23167 19437
rect 23109 19397 23121 19431
rect 23155 19428 23167 19431
rect 23842 19428 23848 19440
rect 23155 19400 23848 19428
rect 23155 19397 23167 19400
rect 23109 19391 23167 19397
rect 23842 19388 23848 19400
rect 23900 19388 23906 19440
rect 26326 19388 26332 19440
rect 26384 19428 26390 19440
rect 28537 19431 28595 19437
rect 28537 19428 28549 19431
rect 26384 19400 28549 19428
rect 26384 19388 26390 19400
rect 28537 19397 28549 19400
rect 28583 19397 28595 19431
rect 28537 19391 28595 19397
rect 29086 19388 29092 19440
rect 29144 19388 29150 19440
rect 31726 19428 31754 19468
rect 32306 19428 32312 19440
rect 31726 19400 32312 19428
rect 32306 19388 32312 19400
rect 32364 19388 32370 19440
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18966 19360 18972 19372
rect 18288 19332 18972 19360
rect 18288 19320 18294 19332
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19116 19332 19257 19360
rect 19116 19320 19122 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 22738 19320 22744 19372
rect 22796 19360 22802 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 22796 19332 24041 19360
rect 22796 19320 22802 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24118 19320 24124 19372
rect 24176 19320 24182 19372
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19329 25007 19363
rect 24949 19323 25007 19329
rect 17880 19264 18000 19292
rect 16482 19224 16488 19236
rect 15948 19196 16488 19224
rect 15841 19187 15899 19193
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 16666 19184 16672 19236
rect 16724 19224 16730 19236
rect 17494 19224 17500 19236
rect 16724 19196 17500 19224
rect 16724 19184 16730 19196
rect 17494 19184 17500 19196
rect 17552 19184 17558 19236
rect 14292 19128 14504 19156
rect 14001 19119 14059 19125
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 15197 19159 15255 19165
rect 15197 19156 15209 19159
rect 15160 19128 15209 19156
rect 15160 19116 15166 19128
rect 15197 19125 15209 19128
rect 15243 19156 15255 19159
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 15243 19128 15393 19156
rect 15243 19125 15255 19128
rect 15197 19119 15255 19125
rect 15381 19125 15393 19128
rect 15427 19156 15439 19159
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15427 19128 16037 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 16025 19125 16037 19128
rect 16071 19156 16083 19159
rect 16206 19156 16212 19168
rect 16071 19128 16212 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 16206 19116 16212 19128
rect 16264 19116 16270 19168
rect 17218 19116 17224 19168
rect 17276 19116 17282 19168
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 17678 19156 17684 19168
rect 17635 19128 17684 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 17972 19156 18000 19264
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 18196 19264 18429 19292
rect 18196 19252 18202 19264
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 22646 19292 22652 19304
rect 20680 19264 22652 19292
rect 20680 19252 20686 19264
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24854 19292 24860 19304
rect 24351 19264 24860 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 18046 19184 18052 19236
rect 18104 19224 18110 19236
rect 19720 19224 19748 19252
rect 18104 19196 19748 19224
rect 18104 19184 18110 19196
rect 22002 19184 22008 19236
rect 22060 19184 22066 19236
rect 22094 19184 22100 19236
rect 22152 19224 22158 19236
rect 23293 19227 23351 19233
rect 23293 19224 23305 19227
rect 22152 19196 23305 19224
rect 22152 19184 22158 19196
rect 23293 19193 23305 19196
rect 23339 19224 23351 19227
rect 24964 19224 24992 19323
rect 26510 19320 26516 19372
rect 26568 19360 26574 19372
rect 27154 19360 27160 19372
rect 26568 19332 27160 19360
rect 26568 19320 26574 19332
rect 27154 19320 27160 19332
rect 27212 19360 27218 19372
rect 27249 19363 27307 19369
rect 27249 19360 27261 19363
rect 27212 19332 27261 19360
rect 27212 19320 27218 19332
rect 27249 19329 27261 19332
rect 27295 19360 27307 19363
rect 27706 19360 27712 19372
rect 27295 19332 27712 19360
rect 27295 19329 27307 19332
rect 27249 19323 27307 19329
rect 27706 19320 27712 19332
rect 27764 19320 27770 19372
rect 30650 19320 30656 19372
rect 30708 19320 30714 19372
rect 25774 19252 25780 19304
rect 25832 19292 25838 19304
rect 27890 19292 27896 19304
rect 25832 19264 27896 19292
rect 25832 19252 25838 19264
rect 27890 19252 27896 19264
rect 27948 19292 27954 19304
rect 28261 19295 28319 19301
rect 28261 19292 28273 19295
rect 27948 19264 28273 19292
rect 27948 19252 27954 19264
rect 28261 19261 28273 19264
rect 28307 19261 28319 19295
rect 28261 19255 28319 19261
rect 25314 19224 25320 19236
rect 23339 19196 23704 19224
rect 23339 19193 23351 19196
rect 23293 19187 23351 19193
rect 17911 19128 18000 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 18782 19116 18788 19168
rect 18840 19156 18846 19168
rect 19968 19159 20026 19165
rect 19968 19156 19980 19159
rect 18840 19128 19980 19156
rect 18840 19116 18846 19128
rect 19968 19125 19980 19128
rect 20014 19156 20026 19159
rect 20990 19156 20996 19168
rect 20014 19128 20996 19156
rect 20014 19125 20026 19128
rect 19968 19119 20026 19125
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 21082 19116 21088 19168
rect 21140 19156 21146 19168
rect 22922 19156 22928 19168
rect 21140 19128 22928 19156
rect 21140 19116 21146 19128
rect 22922 19116 22928 19128
rect 22980 19116 22986 19168
rect 23676 19156 23704 19196
rect 23952 19196 25320 19224
rect 23952 19156 23980 19196
rect 25314 19184 25320 19196
rect 25372 19184 25378 19236
rect 23676 19128 23980 19156
rect 27798 19116 27804 19168
rect 27856 19156 27862 19168
rect 27985 19159 28043 19165
rect 27985 19156 27997 19159
rect 27856 19128 27997 19156
rect 27856 19116 27862 19128
rect 27985 19125 27997 19128
rect 28031 19156 28043 19159
rect 28350 19156 28356 19168
rect 28031 19128 28356 19156
rect 28031 19125 28043 19128
rect 27985 19119 28043 19125
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 30006 19156 30012 19168
rect 28684 19128 30012 19156
rect 28684 19116 28690 19128
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 30282 19116 30288 19168
rect 30340 19156 30346 19168
rect 30929 19159 30987 19165
rect 30929 19156 30941 19159
rect 30340 19128 30941 19156
rect 30340 19116 30346 19128
rect 30929 19125 30941 19128
rect 30975 19125 30987 19159
rect 30929 19119 30987 19125
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 5350 18952 5356 18964
rect 4028 18924 5356 18952
rect 4028 18912 4034 18924
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 7088 18955 7146 18961
rect 7088 18921 7100 18955
rect 7134 18952 7146 18955
rect 7558 18952 7564 18964
rect 7134 18924 7564 18952
rect 7134 18921 7146 18924
rect 7088 18915 7146 18921
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 9401 18955 9459 18961
rect 9401 18952 9413 18955
rect 7892 18924 9413 18952
rect 7892 18912 7898 18924
rect 9401 18921 9413 18924
rect 9447 18921 9459 18955
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 9401 18915 9459 18921
rect 9508 18924 11069 18952
rect 8110 18844 8116 18896
rect 8168 18884 8174 18896
rect 9508 18884 9536 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 11606 18912 11612 18964
rect 11664 18912 11670 18964
rect 14826 18952 14832 18964
rect 11808 18924 14832 18952
rect 8168 18856 9536 18884
rect 8168 18844 8174 18856
rect 10502 18844 10508 18896
rect 10560 18844 10566 18896
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1452 18788 2053 18816
rect 1452 18776 1458 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 2041 18779 2099 18785
rect 4632 18788 6837 18816
rect 4632 18760 4660 18788
rect 6825 18785 6837 18788
rect 6871 18816 6883 18819
rect 8478 18816 8484 18828
rect 6871 18788 8484 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 9030 18816 9036 18828
rect 8812 18788 9036 18816
rect 8812 18776 8818 18788
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 10042 18776 10048 18828
rect 10100 18776 10106 18828
rect 11808 18816 11836 18924
rect 14826 18912 14832 18924
rect 14884 18912 14890 18964
rect 22002 18952 22008 18964
rect 15120 18924 22008 18952
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 14366 18884 14372 18896
rect 12400 18856 14372 18884
rect 12400 18844 12406 18856
rect 14366 18844 14372 18856
rect 14424 18844 14430 18896
rect 10152 18788 11836 18816
rect 10152 18760 10180 18788
rect 12250 18776 12256 18828
rect 12308 18776 12314 18828
rect 13538 18776 13544 18828
rect 13596 18776 13602 18828
rect 13722 18776 13728 18828
rect 13780 18816 13786 18828
rect 15010 18816 15016 18828
rect 13780 18788 15016 18816
rect 13780 18776 13786 18788
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 4522 18748 4528 18760
rect 1811 18720 4528 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18748 9827 18751
rect 10134 18748 10140 18760
rect 9815 18720 10140 18748
rect 9815 18717 9827 18720
rect 9769 18711 9827 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 11848 18720 12817 18748
rect 11848 18708 11854 18720
rect 12805 18717 12817 18720
rect 12851 18748 12863 18751
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 12851 18720 14197 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 14185 18717 14197 18720
rect 14231 18748 14243 18751
rect 14918 18748 14924 18760
rect 14231 18720 14924 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 3896 18652 4752 18680
rect 3896 18624 3924 18652
rect 3605 18615 3663 18621
rect 3605 18581 3617 18615
rect 3651 18612 3663 18615
rect 3878 18612 3884 18624
rect 3651 18584 3884 18612
rect 3651 18581 3663 18584
rect 3605 18575 3663 18581
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 3970 18572 3976 18624
rect 4028 18572 4034 18624
rect 4724 18612 4752 18652
rect 4798 18640 4804 18692
rect 4856 18680 4862 18692
rect 4893 18683 4951 18689
rect 4893 18680 4905 18683
rect 4856 18652 4905 18680
rect 4856 18640 4862 18652
rect 4893 18649 4905 18652
rect 4939 18649 4951 18683
rect 8754 18680 8760 18692
rect 4893 18643 4951 18649
rect 5276 18652 5382 18680
rect 6196 18652 7590 18680
rect 8404 18652 8760 18680
rect 5276 18612 5304 18652
rect 6196 18624 6224 18652
rect 6178 18612 6184 18624
rect 4724 18584 6184 18612
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 6362 18572 6368 18624
rect 6420 18612 6426 18624
rect 8404 18612 8432 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 9950 18680 9956 18692
rect 8864 18652 9956 18680
rect 6420 18584 8432 18612
rect 6420 18572 6426 18584
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 8864 18612 8892 18652
rect 9950 18640 9956 18652
rect 10008 18640 10014 18692
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10965 18683 11023 18689
rect 10965 18680 10977 18683
rect 10284 18652 10977 18680
rect 10284 18640 10290 18652
rect 10965 18649 10977 18652
rect 11011 18680 11023 18683
rect 14553 18683 14611 18689
rect 11011 18652 13952 18680
rect 11011 18649 11023 18652
rect 10965 18643 11023 18649
rect 8628 18584 8892 18612
rect 9125 18615 9183 18621
rect 8628 18572 8634 18584
rect 9125 18581 9137 18615
rect 9171 18612 9183 18615
rect 9861 18615 9919 18621
rect 9861 18612 9873 18615
rect 9171 18584 9873 18612
rect 9171 18581 9183 18584
rect 9125 18575 9183 18581
rect 9861 18581 9873 18584
rect 9907 18612 9919 18615
rect 10410 18612 10416 18624
rect 9907 18584 10416 18612
rect 9907 18581 9919 18584
rect 9861 18575 9919 18581
rect 10410 18572 10416 18584
rect 10468 18572 10474 18624
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11388 18584 11989 18612
rect 11388 18572 11394 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12069 18615 12127 18621
rect 12069 18581 12081 18615
rect 12115 18612 12127 18615
rect 12986 18612 12992 18624
rect 12115 18584 12992 18612
rect 12115 18581 12127 18584
rect 12069 18575 12127 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 13722 18612 13728 18624
rect 13320 18584 13728 18612
rect 13320 18572 13326 18584
rect 13722 18572 13728 18584
rect 13780 18612 13786 18624
rect 13817 18615 13875 18621
rect 13817 18612 13829 18615
rect 13780 18584 13829 18612
rect 13780 18572 13786 18584
rect 13817 18581 13829 18584
rect 13863 18581 13875 18615
rect 13924 18612 13952 18652
rect 14553 18649 14565 18683
rect 14599 18680 14611 18683
rect 15120 18680 15148 18924
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22646 18912 22652 18964
rect 22704 18952 22710 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22704 18924 22937 18952
rect 22704 18912 22710 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23382 18912 23388 18964
rect 23440 18912 23446 18964
rect 23842 18912 23848 18964
rect 23900 18952 23906 18964
rect 24026 18952 24032 18964
rect 23900 18924 24032 18952
rect 23900 18912 23906 18924
rect 24026 18912 24032 18924
rect 24084 18952 24090 18964
rect 25130 18952 25136 18964
rect 24084 18924 25136 18952
rect 24084 18912 24090 18924
rect 25130 18912 25136 18924
rect 25188 18912 25194 18964
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 27157 18955 27215 18961
rect 27157 18952 27169 18955
rect 25740 18924 27169 18952
rect 25740 18912 25746 18924
rect 27157 18921 27169 18924
rect 27203 18921 27215 18955
rect 27157 18915 27215 18921
rect 29086 18912 29092 18964
rect 29144 18952 29150 18964
rect 30282 18952 30288 18964
rect 29144 18924 30288 18952
rect 29144 18912 29150 18924
rect 30282 18912 30288 18924
rect 30340 18952 30346 18964
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 30340 18924 30757 18952
rect 30340 18912 30346 18924
rect 30745 18921 30757 18924
rect 30791 18921 30803 18955
rect 30745 18915 30803 18921
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 18141 18887 18199 18893
rect 16540 18856 17632 18884
rect 16540 18844 16546 18856
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 15243 18788 16712 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 16684 18748 16712 18788
rect 17494 18776 17500 18828
rect 17552 18776 17558 18828
rect 17604 18816 17632 18856
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 18322 18884 18328 18896
rect 18187 18856 18328 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 18322 18844 18328 18856
rect 18380 18844 18386 18896
rect 20162 18844 20168 18896
rect 20220 18884 20226 18896
rect 21082 18884 21088 18896
rect 20220 18856 21088 18884
rect 20220 18844 20226 18856
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 26694 18844 26700 18896
rect 26752 18884 26758 18896
rect 32674 18884 32680 18896
rect 26752 18856 32680 18884
rect 26752 18844 26758 18856
rect 32674 18844 32680 18856
rect 32732 18844 32738 18896
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 17604 18788 18705 18816
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 19760 18788 20361 18816
rect 19760 18776 19766 18788
rect 20349 18785 20361 18788
rect 20395 18816 20407 18819
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20395 18788 21189 18816
rect 20395 18785 20407 18788
rect 20349 18779 20407 18785
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 22002 18776 22008 18828
rect 22060 18816 22066 18828
rect 22060 18788 23520 18816
rect 22060 18776 22066 18788
rect 16850 18748 16856 18760
rect 16684 18720 16856 18748
rect 16850 18708 16856 18720
rect 16908 18748 16914 18760
rect 17126 18748 17132 18760
rect 16908 18720 17132 18748
rect 16908 18708 16914 18720
rect 17126 18708 17132 18720
rect 17184 18748 17190 18760
rect 18046 18748 18052 18760
rect 17184 18720 18052 18748
rect 17184 18708 17190 18720
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 18782 18748 18788 18760
rect 18564 18720 18788 18748
rect 18564 18708 18570 18720
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19659 18720 20852 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 14599 18652 15148 18680
rect 14599 18649 14611 18652
rect 14553 18643 14611 18649
rect 15470 18640 15476 18692
rect 15528 18689 15534 18692
rect 15528 18680 15538 18689
rect 15528 18652 15884 18680
rect 15528 18643 15538 18652
rect 15528 18640 15534 18643
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 13924 18584 14657 18612
rect 13817 18575 13875 18581
rect 14645 18581 14657 18584
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 14921 18615 14979 18621
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15010 18612 15016 18624
rect 14967 18584 15016 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15856 18612 15884 18652
rect 16206 18640 16212 18692
rect 16264 18640 16270 18692
rect 20070 18680 20076 18692
rect 16776 18652 20076 18680
rect 16390 18612 16396 18624
rect 15856 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18612 16454 18624
rect 16776 18612 16804 18652
rect 20070 18640 20076 18652
rect 20128 18640 20134 18692
rect 16448 18584 16804 18612
rect 16448 18572 16454 18584
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 18601 18615 18659 18621
rect 18601 18581 18613 18615
rect 18647 18612 18659 18615
rect 18690 18612 18696 18624
rect 18647 18584 18696 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18612 19395 18615
rect 20254 18612 20260 18624
rect 19383 18584 20260 18612
rect 19383 18581 19395 18584
rect 19337 18575 19395 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20824 18612 20852 18720
rect 20898 18640 20904 18692
rect 20956 18640 20962 18692
rect 23492 18680 23520 18788
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 23716 18788 24593 18816
rect 23716 18776 23722 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25774 18816 25780 18828
rect 25455 18788 25780 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 26142 18776 26148 18828
rect 26200 18816 26206 18828
rect 28718 18816 28724 18828
rect 26200 18788 28724 18816
rect 26200 18776 26206 18788
rect 28718 18776 28724 18788
rect 28776 18776 28782 18828
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 30285 18819 30343 18825
rect 30285 18785 30297 18819
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 26786 18708 26792 18760
rect 26844 18748 26850 18760
rect 27154 18748 27160 18760
rect 26844 18720 27160 18748
rect 26844 18708 26850 18720
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 27614 18708 27620 18760
rect 27672 18708 27678 18760
rect 27893 18751 27951 18757
rect 27893 18717 27905 18751
rect 27939 18748 27951 18751
rect 28902 18748 28908 18760
rect 27939 18720 28908 18748
rect 27939 18717 27951 18720
rect 27893 18711 27951 18717
rect 28902 18708 28908 18720
rect 28960 18708 28966 18760
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 30300 18748 30328 18779
rect 29880 18720 30328 18748
rect 29880 18708 29886 18720
rect 25685 18683 25743 18689
rect 22678 18652 22784 18680
rect 23492 18652 25636 18680
rect 22094 18612 22100 18624
rect 20824 18584 22100 18612
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 22462 18572 22468 18624
rect 22520 18612 22526 18624
rect 22756 18612 22784 18652
rect 24026 18612 24032 18624
rect 22520 18584 24032 18612
rect 22520 18572 22526 18584
rect 24026 18572 24032 18584
rect 24084 18572 24090 18624
rect 24210 18572 24216 18624
rect 24268 18572 24274 18624
rect 25608 18612 25636 18652
rect 25685 18649 25697 18683
rect 25731 18680 25743 18683
rect 25958 18680 25964 18692
rect 25731 18652 25964 18680
rect 25731 18649 25743 18652
rect 25685 18643 25743 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 30742 18680 30748 18692
rect 27080 18652 30748 18680
rect 27080 18612 27108 18652
rect 30742 18640 30748 18652
rect 30800 18640 30806 18692
rect 25608 18584 27108 18612
rect 29730 18572 29736 18624
rect 29788 18572 29794 18624
rect 30098 18572 30104 18624
rect 30156 18572 30162 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 14642 18408 14648 18420
rect 4028 18380 14648 18408
rect 4028 18368 4034 18380
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 15013 18411 15071 18417
rect 15013 18377 15025 18411
rect 15059 18408 15071 18411
rect 15102 18408 15108 18420
rect 15059 18380 15108 18408
rect 15059 18377 15071 18380
rect 15013 18371 15071 18377
rect 15102 18368 15108 18380
rect 15160 18368 15166 18420
rect 16482 18368 16488 18420
rect 16540 18368 16546 18420
rect 17313 18411 17371 18417
rect 17313 18377 17325 18411
rect 17359 18408 17371 18411
rect 20717 18411 20775 18417
rect 20717 18408 20729 18411
rect 17359 18380 20729 18408
rect 17359 18377 17371 18380
rect 17313 18371 17371 18377
rect 20717 18377 20729 18380
rect 20763 18377 20775 18411
rect 20717 18371 20775 18377
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 21048 18380 24869 18408
rect 21048 18368 21054 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 26786 18368 26792 18420
rect 26844 18368 26850 18420
rect 27157 18411 27215 18417
rect 27157 18377 27169 18411
rect 27203 18408 27215 18411
rect 30098 18408 30104 18420
rect 27203 18380 30104 18408
rect 27203 18377 27215 18380
rect 27157 18371 27215 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30834 18368 30840 18420
rect 30892 18408 30898 18420
rect 33318 18408 33324 18420
rect 30892 18380 33324 18408
rect 30892 18368 30898 18380
rect 33318 18368 33324 18380
rect 33376 18368 33382 18420
rect 1780 18312 2774 18340
rect 1780 18281 1808 18312
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 2746 18136 2774 18312
rect 4430 18300 4436 18352
rect 4488 18300 4494 18352
rect 7190 18340 7196 18352
rect 5460 18312 7196 18340
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 5460 18272 5488 18312
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 9766 18300 9772 18352
rect 9824 18300 9830 18352
rect 13998 18340 14004 18352
rect 10980 18312 14004 18340
rect 3651 18244 5488 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 6270 18272 6276 18284
rect 5767 18244 6276 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 6270 18232 6276 18244
rect 6328 18232 6334 18284
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 6914 18272 6920 18284
rect 6779 18244 6920 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 5350 18164 5356 18216
rect 5408 18204 5414 18216
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 5408 18176 5825 18204
rect 5408 18164 5414 18176
rect 5813 18173 5825 18176
rect 5859 18173 5871 18207
rect 5813 18167 5871 18173
rect 5994 18164 6000 18216
rect 6052 18204 6058 18216
rect 7009 18207 7067 18213
rect 7009 18204 7021 18207
rect 6052 18176 7021 18204
rect 6052 18164 6058 18176
rect 7009 18173 7021 18176
rect 7055 18173 7067 18207
rect 7009 18167 7067 18173
rect 7374 18136 7380 18148
rect 2746 18108 7380 18136
rect 7374 18096 7380 18108
rect 7432 18096 7438 18148
rect 8496 18136 8524 18235
rect 10502 18232 10508 18284
rect 10560 18272 10566 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10560 18244 10793 18272
rect 10560 18232 10566 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8628 18176 9229 18204
rect 8628 18164 8634 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9582 18164 9588 18216
rect 9640 18204 9646 18216
rect 10980 18213 11008 18312
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 14461 18343 14519 18349
rect 14461 18309 14473 18343
rect 14507 18340 14519 18343
rect 14550 18340 14556 18352
rect 14507 18312 14556 18340
rect 14507 18309 14519 18312
rect 14461 18303 14519 18309
rect 14550 18300 14556 18312
rect 14608 18300 14614 18352
rect 14826 18300 14832 18352
rect 14884 18340 14890 18352
rect 18141 18343 18199 18349
rect 14884 18312 17540 18340
rect 14884 18300 14890 18312
rect 11882 18232 11888 18284
rect 11940 18272 11946 18284
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 11940 18244 12357 18272
rect 11940 18232 11946 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18272 12495 18275
rect 12618 18272 12624 18284
rect 12483 18244 12624 18272
rect 12483 18241 12495 18244
rect 12437 18235 12495 18241
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13538 18272 13544 18284
rect 13044 18244 13544 18272
rect 13044 18232 13050 18244
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 14918 18272 14924 18284
rect 13679 18244 14924 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 14918 18232 14924 18244
rect 14976 18232 14982 18284
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 15068 18244 15393 18272
rect 15068 18232 15074 18244
rect 15381 18241 15393 18244
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15562 18232 15568 18284
rect 15620 18272 15626 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 15620 18244 17233 18272
rect 15620 18232 15626 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 9640 18176 10885 18204
rect 9640 18164 9646 18176
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 12529 18207 12587 18213
rect 12529 18204 12541 18207
rect 12308 18176 12541 18204
rect 12308 18164 12314 18176
rect 12529 18173 12541 18176
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16942 18204 16948 18216
rect 15703 18176 16948 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 9122 18136 9128 18148
rect 8496 18108 9128 18136
rect 9122 18096 9128 18108
rect 9180 18136 9186 18148
rect 9861 18139 9919 18145
rect 9861 18136 9873 18139
rect 9180 18108 9873 18136
rect 9180 18096 9186 18108
rect 9861 18105 9873 18108
rect 9907 18136 9919 18139
rect 11606 18136 11612 18148
rect 9907 18108 11612 18136
rect 9907 18105 9919 18108
rect 9861 18099 9919 18105
rect 11606 18096 11612 18108
rect 11664 18136 11670 18148
rect 11790 18136 11796 18148
rect 11664 18108 11796 18136
rect 11664 18096 11670 18108
rect 11790 18096 11796 18108
rect 11848 18096 11854 18148
rect 11900 18108 12434 18136
rect 5261 18071 5319 18077
rect 5261 18037 5273 18071
rect 5307 18068 5319 18071
rect 6822 18068 6828 18080
rect 5307 18040 6828 18068
rect 5307 18037 5319 18040
rect 5261 18031 5319 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 10226 18068 10232 18080
rect 6972 18040 10232 18068
rect 6972 18028 6978 18040
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 10413 18071 10471 18077
rect 10413 18037 10425 18071
rect 10459 18068 10471 18071
rect 11900 18068 11928 18108
rect 10459 18040 11928 18068
rect 11977 18071 12035 18077
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12158 18068 12164 18080
rect 12023 18040 12164 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12406 18068 12434 18108
rect 12710 18096 12716 18148
rect 12768 18136 12774 18148
rect 13262 18136 13268 18148
rect 12768 18108 13268 18136
rect 12768 18096 12774 18108
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 15488 18136 15516 18167
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17034 18164 17040 18216
rect 17092 18204 17098 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 17092 18176 17417 18204
rect 17092 18164 17098 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17512 18204 17540 18312
rect 18141 18309 18153 18343
rect 18187 18340 18199 18343
rect 20162 18340 20168 18352
rect 18187 18312 20168 18340
rect 18187 18309 18199 18312
rect 18141 18303 18199 18309
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 21085 18343 21143 18349
rect 21085 18309 21097 18343
rect 21131 18340 21143 18343
rect 22557 18343 22615 18349
rect 22557 18340 22569 18343
rect 21131 18312 22569 18340
rect 21131 18309 21143 18312
rect 21085 18303 21143 18309
rect 22557 18309 22569 18312
rect 22603 18340 22615 18343
rect 22830 18340 22836 18352
rect 22603 18312 22836 18340
rect 22603 18309 22615 18312
rect 22557 18303 22615 18309
rect 17586 18232 17592 18284
rect 17644 18272 17650 18284
rect 19426 18272 19432 18284
rect 17644 18244 19432 18272
rect 17644 18232 17650 18244
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 20254 18272 20260 18284
rect 19935 18244 20260 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 20254 18232 20260 18244
rect 20312 18272 20318 18284
rect 20530 18272 20536 18284
rect 20312 18244 20536 18272
rect 20312 18232 20318 18244
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 17512 18176 18337 18204
rect 17405 18167 17463 18173
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 18325 18167 18383 18173
rect 18877 18207 18935 18213
rect 18877 18173 18889 18207
rect 18923 18204 18935 18207
rect 19610 18204 19616 18216
rect 18923 18176 19616 18204
rect 18923 18173 18935 18176
rect 18877 18167 18935 18173
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 19978 18164 19984 18216
rect 20036 18164 20042 18216
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 19521 18139 19579 18145
rect 19521 18136 19533 18139
rect 15488 18108 19533 18136
rect 19521 18105 19533 18108
rect 19567 18105 19579 18139
rect 19521 18099 19579 18105
rect 20990 18096 20996 18148
rect 21048 18136 21054 18148
rect 21100 18136 21128 18303
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 24026 18300 24032 18352
rect 24084 18300 24090 18352
rect 25314 18300 25320 18352
rect 25372 18300 25378 18352
rect 26050 18300 26056 18352
rect 26108 18300 26114 18352
rect 28353 18343 28411 18349
rect 28353 18309 28365 18343
rect 28399 18340 28411 18343
rect 28626 18340 28632 18352
rect 28399 18312 28632 18340
rect 28399 18309 28411 18312
rect 28353 18303 28411 18309
rect 28626 18300 28632 18312
rect 28684 18300 28690 18352
rect 29086 18300 29092 18352
rect 29144 18300 29150 18352
rect 21174 18232 21180 18284
rect 21232 18232 21238 18284
rect 25332 18272 25360 18300
rect 26513 18275 26571 18281
rect 26513 18272 26525 18275
rect 25332 18244 26525 18272
rect 26513 18241 26525 18244
rect 26559 18241 26571 18275
rect 26513 18235 26571 18241
rect 27798 18232 27804 18284
rect 27856 18272 27862 18284
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 27856 18244 28089 18272
rect 27856 18232 27862 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 30650 18232 30656 18284
rect 30708 18272 30714 18284
rect 41598 18272 41604 18284
rect 30708 18244 31432 18272
rect 30708 18232 30714 18244
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18173 21419 18207
rect 21361 18167 21419 18173
rect 21048 18108 21128 18136
rect 21048 18096 21054 18108
rect 12802 18068 12808 18080
rect 12406 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 16022 18028 16028 18080
rect 16080 18028 16086 18080
rect 16206 18028 16212 18080
rect 16264 18028 16270 18080
rect 16853 18071 16911 18077
rect 16853 18037 16865 18071
rect 16899 18068 16911 18071
rect 17678 18068 17684 18080
rect 16899 18040 17684 18068
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 20622 18028 20628 18080
rect 20680 18068 20686 18080
rect 21376 18068 21404 18167
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21968 18176 22017 18204
rect 21968 18164 21974 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 23109 18207 23167 18213
rect 23109 18173 23121 18207
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 26234 18204 26240 18216
rect 23431 18176 26240 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 20680 18040 21404 18068
rect 20680 18028 20686 18040
rect 21818 18028 21824 18080
rect 21876 18068 21882 18080
rect 22462 18068 22468 18080
rect 21876 18040 22468 18068
rect 21876 18028 21882 18040
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 23124 18068 23152 18167
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 27120 18176 30328 18204
rect 27120 18164 27126 18176
rect 30300 18145 30328 18176
rect 30742 18164 30748 18216
rect 30800 18164 30806 18216
rect 30834 18164 30840 18216
rect 30892 18164 30898 18216
rect 31404 18213 31432 18244
rect 35268 18244 41604 18272
rect 31389 18207 31447 18213
rect 31389 18173 31401 18207
rect 31435 18204 31447 18207
rect 35268 18204 35296 18244
rect 41598 18232 41604 18244
rect 41656 18232 41662 18284
rect 31435 18176 35296 18204
rect 31435 18173 31447 18176
rect 31389 18167 31447 18173
rect 30285 18139 30343 18145
rect 30285 18105 30297 18139
rect 30331 18105 30343 18139
rect 30285 18099 30343 18105
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 30852 18136 30880 18164
rect 30432 18108 30880 18136
rect 30432 18096 30438 18108
rect 24670 18068 24676 18080
rect 23124 18040 24676 18068
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 27338 18028 27344 18080
rect 27396 18068 27402 18080
rect 29822 18068 29828 18080
rect 27396 18040 29828 18068
rect 27396 18028 27402 18040
rect 29822 18028 29828 18040
rect 29880 18028 29886 18080
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 30800 18040 31585 18068
rect 30800 18028 30806 18040
rect 31573 18037 31585 18040
rect 31619 18068 31631 18071
rect 41414 18068 41420 18080
rect 31619 18040 41420 18068
rect 31619 18037 31631 18040
rect 31573 18031 31631 18037
rect 41414 18028 41420 18040
rect 41472 18028 41478 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 3602 17824 3608 17876
rect 3660 17824 3666 17876
rect 3878 17824 3884 17876
rect 3936 17824 3942 17876
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 6641 17867 6699 17873
rect 6641 17864 6653 17867
rect 4856 17836 6653 17864
rect 4856 17824 4862 17836
rect 6641 17833 6653 17836
rect 6687 17833 6699 17867
rect 6641 17827 6699 17833
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7708 17836 7849 17864
rect 7708 17824 7714 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 10376 17836 10609 17864
rect 10376 17824 10382 17836
rect 10597 17833 10609 17836
rect 10643 17833 10655 17867
rect 10597 17827 10655 17833
rect 11606 17824 11612 17876
rect 11664 17824 11670 17876
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13412 17836 13737 17864
rect 13412 17824 13418 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 14458 17824 14464 17876
rect 14516 17824 14522 17876
rect 17126 17864 17132 17876
rect 16316 17836 17132 17864
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 4433 17799 4491 17805
rect 4433 17796 4445 17799
rect 1912 17768 4445 17796
rect 1912 17756 1918 17768
rect 4433 17765 4445 17768
rect 4479 17765 4491 17799
rect 4433 17759 4491 17765
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 7984 17768 11284 17796
rect 7984 17756 7990 17768
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 1780 17700 7389 17728
rect 1780 17669 1808 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 7892 17700 8309 17728
rect 7892 17688 7898 17700
rect 8297 17697 8309 17700
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4614 17660 4620 17672
rect 4212 17632 4620 17660
rect 4212 17620 4218 17632
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4672 17632 4905 17660
rect 4672 17620 4678 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 7098 17620 7104 17672
rect 7156 17660 7162 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7156 17632 8217 17660
rect 7156 17620 7162 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8404 17660 8432 17691
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9456 17700 9873 17728
rect 9456 17688 9462 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10008 17700 11161 17728
rect 10008 17688 10014 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11256 17728 11284 17768
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 14366 17796 14372 17808
rect 13320 17768 14372 17796
rect 13320 17756 13326 17768
rect 14366 17756 14372 17768
rect 14424 17756 14430 17808
rect 16114 17728 16120 17740
rect 11256 17700 16120 17728
rect 11149 17691 11207 17697
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 16316 17737 16344 17836
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 17310 17824 17316 17876
rect 17368 17864 17374 17876
rect 19659 17867 19717 17873
rect 19659 17864 19671 17867
rect 17368 17836 19671 17864
rect 17368 17824 17374 17836
rect 19659 17833 19671 17836
rect 19705 17833 19717 17867
rect 19659 17827 19717 17833
rect 21818 17824 21824 17876
rect 21876 17824 21882 17876
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 27522 17864 27528 17876
rect 21968 17836 27528 17864
rect 21968 17824 21974 17836
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 28626 17824 28632 17876
rect 28684 17864 28690 17876
rect 28810 17864 28816 17876
rect 28684 17836 28816 17864
rect 28684 17824 28690 17836
rect 28810 17824 28816 17836
rect 28868 17824 28874 17876
rect 17586 17756 17592 17808
rect 17644 17796 17650 17808
rect 20717 17799 20775 17805
rect 20717 17796 20729 17799
rect 17644 17768 20729 17796
rect 17644 17756 17650 17768
rect 20717 17765 20729 17768
rect 20763 17765 20775 17799
rect 20717 17759 20775 17765
rect 21082 17756 21088 17808
rect 21140 17796 21146 17808
rect 22002 17796 22008 17808
rect 21140 17768 22008 17796
rect 21140 17756 21146 17768
rect 22002 17756 22008 17768
rect 22060 17756 22066 17808
rect 26234 17756 26240 17808
rect 26292 17796 26298 17808
rect 26605 17799 26663 17805
rect 26605 17796 26617 17799
rect 26292 17768 26617 17796
rect 26292 17756 26298 17768
rect 26605 17765 26617 17768
rect 26651 17765 26663 17799
rect 26605 17759 26663 17765
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 29733 17799 29791 17805
rect 29733 17796 29745 17799
rect 28500 17768 29745 17796
rect 28500 17756 28506 17768
rect 29733 17765 29745 17768
rect 29779 17765 29791 17799
rect 30374 17796 30380 17808
rect 29733 17759 29791 17765
rect 30300 17768 30380 17796
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16942 17728 16948 17740
rect 16623 17700 16948 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 17218 17688 17224 17740
rect 17276 17728 17282 17740
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 17276 17700 19441 17728
rect 17276 17688 17282 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 20404 17700 21281 17728
rect 20404 17688 20410 17700
rect 21269 17697 21281 17700
rect 21315 17728 21327 17731
rect 24578 17728 24584 17740
rect 21315 17700 24584 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 24578 17688 24584 17700
rect 24636 17688 24642 17740
rect 24670 17688 24676 17740
rect 24728 17728 24734 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24728 17700 24869 17728
rect 24728 17688 24734 17700
rect 24857 17697 24869 17700
rect 24903 17728 24915 17731
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 24903 17700 27077 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 27065 17697 27077 17700
rect 27111 17728 27123 17731
rect 27798 17728 27804 17740
rect 27111 17700 27804 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 27798 17688 27804 17700
rect 27856 17688 27862 17740
rect 29178 17728 29184 17740
rect 28460 17700 29184 17728
rect 10226 17660 10232 17672
rect 8205 17623 8263 17629
rect 8312 17632 10232 17660
rect 1210 17552 1216 17604
rect 1268 17592 1274 17604
rect 2501 17595 2559 17601
rect 2501 17592 2513 17595
rect 1268 17564 2513 17592
rect 1268 17552 1274 17564
rect 2501 17561 2513 17564
rect 2547 17561 2559 17595
rect 2501 17555 2559 17561
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17592 4307 17595
rect 4338 17592 4344 17604
rect 4295 17564 4344 17592
rect 4295 17561 4307 17564
rect 4249 17555 4307 17561
rect 4338 17552 4344 17564
rect 4396 17552 4402 17604
rect 5169 17595 5227 17601
rect 5169 17561 5181 17595
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 5184 17524 5212 17555
rect 6178 17552 6184 17604
rect 6236 17552 6242 17604
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 7466 17592 7472 17604
rect 7239 17564 7472 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 7466 17552 7472 17564
rect 7524 17552 7530 17604
rect 7558 17552 7564 17604
rect 7616 17592 7622 17604
rect 8312 17592 8340 17632
rect 10226 17620 10232 17632
rect 10284 17660 10290 17672
rect 10870 17660 10876 17672
rect 10284 17632 10876 17660
rect 10284 17620 10290 17632
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 10962 17620 10968 17672
rect 11020 17620 11026 17672
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 20622 17660 20628 17672
rect 18524 17632 20628 17660
rect 7616 17564 8340 17592
rect 7616 17552 7622 17564
rect 9122 17552 9128 17604
rect 9180 17552 9186 17604
rect 9646 17564 12204 17592
rect 8294 17524 8300 17536
rect 5184 17496 8300 17524
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 9646 17524 9674 17564
rect 8444 17496 9674 17524
rect 8444 17484 8450 17496
rect 10686 17484 10692 17536
rect 10744 17524 10750 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10744 17496 11069 17524
rect 10744 17484 10750 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 12176 17524 12204 17564
rect 12250 17552 12256 17604
rect 12308 17552 12314 17604
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 16206 17592 16212 17604
rect 14415 17564 14872 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 14844 17536 14872 17564
rect 15948 17564 16212 17592
rect 15948 17536 15976 17564
rect 16206 17552 16212 17564
rect 16264 17592 16270 17604
rect 18325 17595 18383 17601
rect 18325 17592 18337 17595
rect 16264 17564 17066 17592
rect 17880 17564 18337 17592
rect 16264 17552 16270 17564
rect 14090 17524 14096 17536
rect 12176 17496 14096 17524
rect 11057 17487 11115 17493
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14826 17484 14832 17536
rect 14884 17484 14890 17536
rect 14918 17484 14924 17536
rect 14976 17524 14982 17536
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 14976 17496 15025 17524
rect 14976 17484 14982 17496
rect 15013 17493 15025 17496
rect 15059 17493 15071 17527
rect 15013 17487 15071 17493
rect 15378 17484 15384 17536
rect 15436 17484 15442 17536
rect 15930 17484 15936 17536
rect 15988 17484 15994 17536
rect 16960 17524 16988 17564
rect 17880 17524 17908 17564
rect 18325 17561 18337 17564
rect 18371 17561 18383 17595
rect 18325 17555 18383 17561
rect 18524 17536 18552 17632
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 21174 17620 21180 17672
rect 21232 17620 21238 17672
rect 22002 17620 22008 17672
rect 22060 17660 22066 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22060 17632 22293 17660
rect 22060 17620 22066 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 24026 17660 24032 17672
rect 23690 17632 24032 17660
rect 22281 17623 22339 17629
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 28460 17646 28488 17700
rect 29178 17688 29184 17700
rect 29236 17688 29242 17740
rect 30190 17688 30196 17740
rect 30248 17688 30254 17740
rect 30300 17737 30328 17768
rect 30374 17756 30380 17768
rect 30432 17756 30438 17808
rect 30285 17731 30343 17737
rect 30285 17697 30297 17731
rect 30331 17697 30343 17731
rect 31481 17731 31539 17737
rect 31481 17728 31493 17731
rect 30285 17691 30343 17697
rect 30392 17700 31493 17728
rect 30392 17660 30420 17700
rect 31481 17697 31493 17700
rect 31527 17697 31539 17731
rect 31481 17691 31539 17697
rect 28828 17632 30420 17660
rect 19610 17552 19616 17604
rect 19668 17592 19674 17604
rect 21085 17595 21143 17601
rect 21085 17592 21097 17595
rect 19668 17564 21097 17592
rect 19668 17552 19674 17564
rect 21085 17561 21097 17564
rect 21131 17561 21143 17595
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 21085 17555 21143 17561
rect 21192 17564 22569 17592
rect 16960 17496 17908 17524
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18506 17524 18512 17536
rect 18095 17496 18512 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 20438 17524 20444 17536
rect 18739 17496 20444 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20622 17484 20628 17536
rect 20680 17524 20686 17536
rect 21192 17524 21220 17564
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 24394 17592 24400 17604
rect 22557 17555 22615 17561
rect 23952 17564 24400 17592
rect 20680 17496 21220 17524
rect 20680 17484 20686 17496
rect 21910 17484 21916 17536
rect 21968 17484 21974 17536
rect 23566 17484 23572 17536
rect 23624 17524 23630 17536
rect 23952 17524 23980 17564
rect 24394 17552 24400 17564
rect 24452 17552 24458 17604
rect 25130 17552 25136 17604
rect 25188 17552 25194 17604
rect 26786 17592 26792 17604
rect 26358 17564 26792 17592
rect 26786 17552 26792 17564
rect 26844 17552 26850 17604
rect 27338 17552 27344 17604
rect 27396 17552 27402 17604
rect 23624 17496 23980 17524
rect 24029 17527 24087 17533
rect 23624 17484 23630 17496
rect 24029 17493 24041 17527
rect 24075 17524 24087 17527
rect 25148 17524 25176 17552
rect 28828 17536 28856 17632
rect 30834 17620 30840 17672
rect 30892 17660 30898 17672
rect 31202 17660 31208 17672
rect 30892 17632 31208 17660
rect 30892 17620 30898 17632
rect 31202 17620 31208 17632
rect 31260 17660 31266 17672
rect 31297 17663 31355 17669
rect 31297 17660 31309 17663
rect 31260 17632 31309 17660
rect 31260 17620 31266 17632
rect 31297 17629 31309 17632
rect 31343 17629 31355 17663
rect 31297 17623 31355 17629
rect 31389 17663 31447 17669
rect 31389 17629 31401 17663
rect 31435 17660 31447 17663
rect 34698 17660 34704 17672
rect 31435 17632 34704 17660
rect 31435 17629 31447 17632
rect 31389 17623 31447 17629
rect 34698 17620 34704 17632
rect 34756 17620 34762 17672
rect 30098 17552 30104 17604
rect 30156 17552 30162 17604
rect 24075 17496 25176 17524
rect 24075 17493 24087 17496
rect 24029 17487 24087 17493
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 27614 17524 27620 17536
rect 25280 17496 27620 17524
rect 25280 17484 25286 17496
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 28810 17484 28816 17536
rect 28868 17484 28874 17536
rect 29178 17484 29184 17536
rect 29236 17484 29242 17536
rect 30926 17484 30932 17536
rect 30984 17484 30990 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 5307 17292 7297 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7432 17292 8033 17320
rect 7432 17280 7438 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 8110 17280 8116 17332
rect 8168 17320 8174 17332
rect 8386 17320 8392 17332
rect 8168 17292 8392 17320
rect 8168 17280 8174 17292
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 8481 17323 8539 17329
rect 8481 17289 8493 17323
rect 8527 17320 8539 17323
rect 9766 17320 9772 17332
rect 8527 17292 9772 17320
rect 8527 17289 8539 17292
rect 8481 17283 8539 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 11241 17323 11299 17329
rect 11241 17320 11253 17323
rect 9916 17292 11253 17320
rect 9916 17280 9922 17292
rect 11241 17289 11253 17292
rect 11287 17320 11299 17323
rect 12066 17320 12072 17332
rect 11287 17292 12072 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12526 17280 12532 17332
rect 12584 17280 12590 17332
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 14148 17292 14197 17320
rect 14148 17280 14154 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 16114 17280 16120 17332
rect 16172 17280 16178 17332
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 22005 17323 22063 17329
rect 22005 17320 22017 17323
rect 17920 17292 22017 17320
rect 17920 17280 17926 17292
rect 22005 17289 22017 17292
rect 22051 17289 22063 17323
rect 22005 17283 22063 17289
rect 22373 17323 22431 17329
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 22830 17320 22836 17332
rect 22419 17292 22836 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 23566 17280 23572 17332
rect 23624 17320 23630 17332
rect 23661 17323 23719 17329
rect 23661 17320 23673 17323
rect 23624 17292 23673 17320
rect 23624 17280 23630 17292
rect 23661 17289 23673 17292
rect 23707 17289 23719 17323
rect 23661 17283 23719 17289
rect 23753 17323 23811 17329
rect 23753 17289 23765 17323
rect 23799 17320 23811 17323
rect 24210 17320 24216 17332
rect 23799 17292 24216 17320
rect 23799 17289 23811 17292
rect 23753 17283 23811 17289
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 28810 17320 28816 17332
rect 24964 17292 28816 17320
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 4982 17252 4988 17264
rect 4663 17224 4988 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 6512 17224 10977 17252
rect 6512 17212 6518 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 12894 17212 12900 17264
rect 12952 17212 12958 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 14016 17224 14749 17252
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 3651 17156 4752 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 4724 17048 4752 17156
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 5721 17187 5779 17193
rect 5721 17153 5733 17187
rect 5767 17184 5779 17187
rect 5767 17156 5948 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 5920 17128 5948 17156
rect 6178 17144 6184 17196
rect 6236 17184 6242 17196
rect 6362 17184 6368 17196
rect 6236 17156 6368 17184
rect 6236 17144 6242 17156
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9582 17184 9588 17196
rect 9088 17156 9588 17184
rect 9088 17144 9094 17156
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 9950 17144 9956 17196
rect 10008 17144 10014 17196
rect 10781 17188 10839 17193
rect 10870 17188 10876 17196
rect 10781 17187 10876 17188
rect 10781 17153 10793 17187
rect 10827 17160 10876 17187
rect 10827 17153 10839 17160
rect 10781 17147 10839 17153
rect 10870 17144 10876 17160
rect 10928 17144 10934 17196
rect 11146 17144 11152 17196
rect 11204 17184 11210 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11204 17156 11805 17184
rect 11204 17144 11210 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 14016 17184 14044 17224
rect 14737 17221 14749 17224
rect 14783 17252 14795 17255
rect 18690 17252 18696 17264
rect 14783 17224 18696 17252
rect 14783 17221 14795 17224
rect 14737 17215 14795 17221
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 20162 17212 20168 17264
rect 20220 17252 20226 17264
rect 21085 17255 21143 17261
rect 21085 17252 21097 17255
rect 20220 17224 21097 17252
rect 20220 17212 20226 17224
rect 21085 17221 21097 17224
rect 21131 17252 21143 17255
rect 21910 17252 21916 17264
rect 21131 17224 21916 17252
rect 21131 17221 21143 17224
rect 21085 17215 21143 17221
rect 21910 17212 21916 17224
rect 21968 17252 21974 17264
rect 24964 17261 24992 17292
rect 28810 17280 28816 17292
rect 28868 17280 28874 17332
rect 30098 17280 30104 17332
rect 30156 17320 30162 17332
rect 30282 17320 30288 17332
rect 30156 17292 30288 17320
rect 30156 17280 30162 17292
rect 30282 17280 30288 17292
rect 30340 17320 30346 17332
rect 30929 17323 30987 17329
rect 30929 17320 30941 17323
rect 30340 17292 30941 17320
rect 30340 17280 30346 17292
rect 30929 17289 30941 17292
rect 30975 17289 30987 17323
rect 30929 17283 30987 17289
rect 22465 17255 22523 17261
rect 22465 17252 22477 17255
rect 21968 17224 22477 17252
rect 21968 17212 21974 17224
rect 22465 17221 22477 17224
rect 22511 17221 22523 17255
rect 22465 17215 22523 17221
rect 24949 17255 25007 17261
rect 24949 17221 24961 17255
rect 24995 17221 25007 17255
rect 26786 17252 26792 17264
rect 26174 17224 26792 17252
rect 24949 17215 25007 17221
rect 26786 17212 26792 17224
rect 26844 17212 26850 17264
rect 30190 17212 30196 17264
rect 30248 17252 30254 17264
rect 30561 17255 30619 17261
rect 30561 17252 30573 17255
rect 30248 17224 30573 17252
rect 30248 17212 30254 17224
rect 30561 17221 30573 17224
rect 30607 17252 30619 17255
rect 30607 17224 31754 17252
rect 30607 17221 30619 17224
rect 30561 17215 30619 17221
rect 11793 17147 11851 17153
rect 13096 17156 14044 17184
rect 5810 17076 5816 17128
rect 5868 17076 5874 17128
rect 5902 17076 5908 17128
rect 5960 17076 5966 17128
rect 7469 17119 7527 17125
rect 6012 17088 6960 17116
rect 6012 17048 6040 17088
rect 4724 17020 6040 17048
rect 6730 17008 6736 17060
rect 6788 17048 6794 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 6788 17020 6837 17048
rect 6788 17008 6794 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6932 17048 6960 17088
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7558 17116 7564 17128
rect 7515 17088 7564 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8754 17116 8760 17128
rect 8711 17088 8760 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 8938 17076 8944 17128
rect 8996 17116 9002 17128
rect 9968 17116 9996 17144
rect 8996 17088 9996 17116
rect 10045 17119 10103 17125
rect 8996 17076 9002 17088
rect 10045 17085 10057 17119
rect 10091 17085 10103 17119
rect 10045 17079 10103 17085
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17116 13047 17119
rect 13096 17116 13124 17156
rect 14090 17144 14096 17196
rect 14148 17144 14154 17196
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 17126 17184 17132 17196
rect 16347 17156 17132 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17218 17144 17224 17196
rect 17276 17144 17282 17196
rect 21818 17184 21824 17196
rect 19550 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 27798 17144 27804 17196
rect 27856 17144 27862 17196
rect 29178 17144 29184 17196
rect 29236 17184 29242 17196
rect 30098 17184 30104 17196
rect 29236 17156 30104 17184
rect 29236 17144 29242 17156
rect 30098 17144 30104 17156
rect 30156 17144 30162 17196
rect 30834 17144 30840 17196
rect 30892 17144 30898 17196
rect 13035 17088 13124 17116
rect 13173 17119 13231 17125
rect 13035 17085 13047 17088
rect 12989 17079 13047 17085
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13354 17116 13360 17128
rect 13219 17088 13360 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 6932 17020 9674 17048
rect 6825 17011 6883 17017
rect 4338 16940 4344 16992
rect 4396 16980 4402 16992
rect 6178 16980 6184 16992
rect 4396 16952 6184 16980
rect 4396 16940 4402 16952
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6549 16983 6607 16989
rect 6549 16949 6561 16983
rect 6595 16980 6607 16983
rect 7466 16980 7472 16992
rect 6595 16952 7472 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 7834 16980 7840 16992
rect 7616 16952 7840 16980
rect 7616 16940 7622 16952
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 9030 16980 9036 16992
rect 8812 16952 9036 16980
rect 8812 16940 8818 16952
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 9646 16980 9674 17020
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 10060 17048 10088 17079
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 15470 17116 15476 17128
rect 14415 17088 15476 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 15838 17076 15844 17128
rect 15896 17116 15902 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 15896 17088 17325 17116
rect 15896 17076 15902 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 18506 17116 18512 17128
rect 18463 17088 18512 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 10318 17048 10324 17060
rect 9824 17020 10324 17048
rect 9824 17008 9830 17020
rect 10318 17008 10324 17020
rect 10376 17008 10382 17060
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 13725 17051 13783 17057
rect 11848 17020 13400 17048
rect 11848 17008 11854 17020
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 9646 16952 11897 16980
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 12434 16980 12440 16992
rect 12124 16952 12440 16980
rect 12124 16940 12130 16952
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 13262 16980 13268 16992
rect 12584 16952 13268 16980
rect 12584 16940 12590 16952
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 13372 16980 13400 17020
rect 13725 17017 13737 17051
rect 13771 17048 13783 17051
rect 15010 17048 15016 17060
rect 13771 17020 15016 17048
rect 13771 17017 13783 17020
rect 13725 17011 13783 17017
rect 15010 17008 15016 17020
rect 15068 17008 15074 17060
rect 16853 17051 16911 17057
rect 16853 17048 16865 17051
rect 15120 17020 16865 17048
rect 15120 16980 15148 17020
rect 16853 17017 16865 17020
rect 16899 17017 16911 17051
rect 16853 17011 16911 17017
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 18156 17048 18184 17079
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 18782 17076 18788 17128
rect 18840 17116 18846 17128
rect 20990 17116 20996 17128
rect 18840 17088 20996 17116
rect 18840 17076 18846 17088
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 21082 17076 21088 17128
rect 21140 17116 21146 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 21140 17088 21189 17116
rect 21140 17076 21146 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17085 21419 17119
rect 21361 17079 21419 17085
rect 20622 17048 20628 17060
rect 17092 17020 18184 17048
rect 19904 17020 20628 17048
rect 17092 17008 17098 17020
rect 13372 16952 15148 16980
rect 15470 16940 15476 16992
rect 15528 16940 15534 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 19904 16989 19932 17020
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 20714 17008 20720 17060
rect 20772 17008 20778 17060
rect 21376 17048 21404 17079
rect 22554 17076 22560 17128
rect 22612 17076 22618 17128
rect 23845 17119 23903 17125
rect 23845 17085 23857 17119
rect 23891 17085 23903 17119
rect 23845 17079 23903 17085
rect 22646 17048 22652 17060
rect 21376 17020 22652 17048
rect 22646 17008 22652 17020
rect 22704 17048 22710 17060
rect 23860 17048 23888 17079
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 26421 17119 26479 17125
rect 26421 17116 26433 17119
rect 24636 17088 26433 17116
rect 24636 17076 24642 17088
rect 26421 17085 26433 17088
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27706 17116 27712 17128
rect 27203 17088 27712 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 27706 17076 27712 17088
rect 27764 17076 27770 17128
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 30374 17116 30380 17128
rect 28123 17088 30380 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 22704 17020 23888 17048
rect 31726 17048 31754 17224
rect 45278 17048 45284 17060
rect 31726 17020 45284 17048
rect 22704 17008 22710 17020
rect 45278 17008 45284 17020
rect 45336 17008 45342 17060
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 17000 16952 19901 16980
rect 17000 16940 17006 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 20070 16940 20076 16992
rect 20128 16980 20134 16992
rect 20349 16983 20407 16989
rect 20349 16980 20361 16983
rect 20128 16952 20361 16980
rect 20128 16940 20134 16952
rect 20349 16949 20361 16952
rect 20395 16980 20407 16983
rect 21082 16980 21088 16992
rect 20395 16952 21088 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21358 16940 21364 16992
rect 21416 16980 21422 16992
rect 22738 16980 22744 16992
rect 21416 16952 22744 16980
rect 21416 16940 21422 16952
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 23290 16940 23296 16992
rect 23348 16940 23354 16992
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 26142 16980 26148 16992
rect 24452 16952 26148 16980
rect 24452 16940 24458 16952
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 29549 16983 29607 16989
rect 29549 16980 29561 16983
rect 27304 16952 29561 16980
rect 27304 16940 27310 16952
rect 29549 16949 29561 16952
rect 29595 16949 29607 16983
rect 29549 16943 29607 16949
rect 29917 16983 29975 16989
rect 29917 16949 29929 16983
rect 29963 16980 29975 16983
rect 30098 16980 30104 16992
rect 29963 16952 30104 16980
rect 29963 16949 29975 16952
rect 29917 16943 29975 16949
rect 30098 16940 30104 16952
rect 30156 16940 30162 16992
rect 30282 16940 30288 16992
rect 30340 16980 30346 16992
rect 48774 16980 48780 16992
rect 30340 16952 48780 16980
rect 30340 16940 30346 16952
rect 48774 16940 48780 16952
rect 48832 16940 48838 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 5718 16736 5724 16788
rect 5776 16776 5782 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5776 16748 6009 16776
rect 5776 16736 5782 16748
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 5997 16739 6055 16745
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 7558 16776 7564 16788
rect 6236 16748 7564 16776
rect 6236 16736 6242 16748
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 7668 16748 7972 16776
rect 7668 16708 7696 16748
rect 3712 16680 7696 16708
rect 7944 16708 7972 16748
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8076 16748 13492 16776
rect 8076 16736 8082 16748
rect 9401 16711 9459 16717
rect 9401 16708 9413 16711
rect 7944 16680 9413 16708
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 3712 16572 3740 16680
rect 9401 16677 9413 16680
rect 9447 16677 9459 16711
rect 9401 16671 9459 16677
rect 9769 16711 9827 16717
rect 9769 16677 9781 16711
rect 9815 16708 9827 16711
rect 10410 16708 10416 16720
rect 9815 16680 10416 16708
rect 9815 16677 9827 16680
rect 9769 16671 9827 16677
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 12894 16708 12900 16720
rect 12308 16680 12900 16708
rect 12308 16668 12314 16680
rect 12894 16668 12900 16680
rect 12952 16668 12958 16720
rect 6730 16600 6736 16652
rect 6788 16640 6794 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 6788 16612 7113 16640
rect 6788 16600 6794 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 7331 16612 7788 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 1811 16544 3740 16572
rect 3973 16575 4031 16581
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 5905 16575 5963 16581
rect 5905 16541 5917 16575
rect 5951 16572 5963 16575
rect 7650 16572 7656 16584
rect 5951 16544 7656 16572
rect 5951 16541 5963 16544
rect 5905 16535 5963 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2501 16467 2559 16473
rect 3988 16436 4016 16535
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7760 16572 7788 16612
rect 7944 16612 8493 16640
rect 7944 16572 7972 16612
rect 8481 16609 8493 16612
rect 8527 16640 8539 16643
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 8527 16612 10701 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 10689 16609 10701 16612
rect 10735 16640 10747 16643
rect 10735 16612 11100 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 7760 16544 7972 16572
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8297 16575 8355 16581
rect 8297 16572 8309 16575
rect 8168 16544 8309 16572
rect 8168 16532 8174 16544
rect 8297 16541 8309 16544
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 10192 16544 10425 16572
rect 10192 16532 10198 16544
rect 10413 16541 10425 16544
rect 10459 16541 10471 16575
rect 11072 16572 11100 16612
rect 11330 16600 11336 16652
rect 11388 16640 11394 16652
rect 13464 16649 13492 16748
rect 14366 16736 14372 16788
rect 14424 16776 14430 16788
rect 18874 16776 18880 16788
rect 14424 16748 18880 16776
rect 14424 16736 14430 16748
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 30926 16776 30932 16788
rect 21232 16748 30932 16776
rect 21232 16736 21238 16748
rect 30926 16736 30932 16748
rect 30984 16736 30990 16788
rect 18506 16708 18512 16720
rect 13648 16680 18512 16708
rect 13648 16649 13676 16680
rect 18506 16668 18512 16680
rect 18564 16668 18570 16720
rect 23566 16708 23572 16720
rect 22664 16680 23572 16708
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 11388 16612 11713 16640
rect 11388 16600 11394 16612
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 11900 16572 11928 16603
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15252 16612 15485 16640
rect 15252 16600 15258 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 16298 16640 16304 16652
rect 15703 16612 16304 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16640 16819 16643
rect 17218 16640 17224 16652
rect 16807 16612 17224 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20346 16640 20352 16652
rect 19751 16612 20352 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 22664 16649 22692 16680
rect 23566 16668 23572 16680
rect 23624 16668 23630 16720
rect 25130 16668 25136 16720
rect 25188 16708 25194 16720
rect 25188 16680 28488 16708
rect 25188 16668 25194 16680
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 20772 16612 22477 16640
rect 20772 16600 20778 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22649 16643 22707 16649
rect 22649 16609 22661 16643
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 22830 16600 22836 16652
rect 22888 16640 22894 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 22888 16612 23765 16640
rect 22888 16600 22894 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23842 16600 23848 16652
rect 23900 16600 23906 16652
rect 25222 16600 25228 16652
rect 25280 16600 25286 16652
rect 25314 16600 25320 16652
rect 25372 16640 25378 16652
rect 25777 16643 25835 16649
rect 25777 16640 25789 16643
rect 25372 16612 25789 16640
rect 25372 16600 25378 16612
rect 25777 16609 25789 16612
rect 25823 16640 25835 16643
rect 25866 16640 25872 16652
rect 25823 16612 25872 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 25866 16600 25872 16612
rect 25924 16600 25930 16652
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27246 16600 27252 16652
rect 27304 16600 27310 16652
rect 28460 16649 28488 16680
rect 28626 16668 28632 16720
rect 28684 16708 28690 16720
rect 30834 16708 30840 16720
rect 28684 16680 30840 16708
rect 28684 16668 28690 16680
rect 30834 16668 30840 16680
rect 30892 16668 30898 16720
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 31294 16640 31300 16652
rect 28491 16612 31300 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 31294 16600 31300 16612
rect 31352 16600 31358 16652
rect 12342 16572 12348 16584
rect 11072 16544 12348 16572
rect 10413 16535 10471 16541
rect 12342 16532 12348 16544
rect 12400 16572 12406 16584
rect 12434 16572 12440 16584
rect 12400 16544 12440 16572
rect 12400 16532 12406 16544
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 14826 16572 14832 16584
rect 14599 16544 14832 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 15378 16532 15384 16584
rect 15436 16532 15442 16584
rect 16574 16532 16580 16584
rect 16632 16572 16638 16584
rect 17310 16572 17316 16584
rect 16632 16544 17316 16572
rect 16632 16532 16638 16544
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16572 18291 16575
rect 18322 16572 18328 16584
rect 18279 16544 18328 16572
rect 18279 16541 18291 16544
rect 18233 16535 18291 16541
rect 5166 16464 5172 16516
rect 5224 16464 5230 16516
rect 7742 16504 7748 16516
rect 5920 16476 7748 16504
rect 5920 16436 5948 16476
rect 7742 16464 7748 16476
rect 7800 16464 7806 16516
rect 9030 16504 9036 16516
rect 7852 16476 9036 16504
rect 3988 16408 5948 16436
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6730 16436 6736 16448
rect 6687 16408 6736 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7852 16445 7880 16476
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 9217 16507 9275 16513
rect 9217 16473 9229 16507
rect 9263 16504 9275 16507
rect 12158 16504 12164 16516
rect 9263 16476 12164 16504
rect 9263 16473 9275 16476
rect 9217 16467 9275 16473
rect 12158 16464 12164 16476
rect 12216 16464 12222 16516
rect 12802 16464 12808 16516
rect 12860 16504 12866 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12860 16476 13369 16504
rect 12860 16464 12866 16476
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 15562 16504 15568 16516
rect 13357 16467 13415 16473
rect 14292 16476 15568 16504
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6972 16408 7021 16436
rect 6972 16396 6978 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7009 16399 7067 16405
rect 7837 16439 7895 16445
rect 7837 16405 7849 16439
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 8754 16436 8760 16448
rect 8251 16408 8760 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 10045 16439 10103 16445
rect 10045 16436 10057 16439
rect 9824 16408 10057 16436
rect 9824 16396 9830 16408
rect 10045 16405 10057 16408
rect 10091 16405 10103 16439
rect 10045 16399 10103 16405
rect 10410 16396 10416 16448
rect 10468 16436 10474 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10468 16408 10517 16436
rect 10468 16396 10474 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 11238 16396 11244 16448
rect 11296 16396 11302 16448
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16436 11667 16439
rect 11698 16436 11704 16448
rect 11655 16408 11704 16436
rect 11655 16405 11667 16408
rect 11609 16399 11667 16405
rect 11698 16396 11704 16408
rect 11756 16436 11762 16448
rect 12253 16439 12311 16445
rect 12253 16436 12265 16439
rect 11756 16408 12265 16436
rect 11756 16396 11762 16408
rect 12253 16405 12265 16408
rect 12299 16405 12311 16439
rect 12253 16399 12311 16405
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16436 13047 16439
rect 14292 16436 14320 16476
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 17604 16504 17632 16535
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 18656 16544 18705 16572
rect 18656 16532 18662 16544
rect 18693 16541 18705 16544
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 21818 16572 21824 16584
rect 20838 16544 21824 16572
rect 21818 16532 21824 16544
rect 21876 16532 21882 16584
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 23290 16572 23296 16584
rect 22419 16544 23296 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 23860 16572 23888 16600
rect 24026 16572 24032 16584
rect 23707 16544 24032 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 24026 16532 24032 16544
rect 24084 16532 24090 16584
rect 25038 16532 25044 16584
rect 25096 16572 25102 16584
rect 25096 16544 26740 16572
rect 25096 16532 25102 16544
rect 17604 16476 19656 16504
rect 13035 16408 14320 16436
rect 13035 16405 13047 16408
rect 12989 16399 13047 16405
rect 14366 16396 14372 16448
rect 14424 16396 14430 16448
rect 15013 16439 15071 16445
rect 15013 16405 15025 16439
rect 15059 16436 15071 16439
rect 16482 16436 16488 16448
rect 15059 16408 16488 16436
rect 15059 16405 15071 16408
rect 15013 16399 15071 16405
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 16666 16396 16672 16448
rect 16724 16436 16730 16448
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 16724 16408 17417 16436
rect 16724 16396 16730 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18049 16439 18107 16445
rect 18049 16405 18061 16439
rect 18095 16436 18107 16439
rect 19518 16436 19524 16448
rect 18095 16408 19524 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 19628 16436 19656 16476
rect 21450 16464 21456 16516
rect 21508 16464 21514 16516
rect 23842 16504 23848 16516
rect 21560 16476 23848 16504
rect 21560 16436 21588 16476
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24176 16476 26648 16504
rect 24176 16464 24182 16476
rect 19628 16408 21588 16436
rect 21634 16396 21640 16448
rect 21692 16436 21698 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21692 16408 22017 16436
rect 21692 16396 21698 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 22520 16408 23213 16436
rect 22520 16396 22526 16408
rect 23201 16405 23213 16408
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 23474 16396 23480 16448
rect 23532 16436 23538 16448
rect 23569 16439 23627 16445
rect 23569 16436 23581 16439
rect 23532 16408 23581 16436
rect 23532 16396 23538 16408
rect 23569 16405 23581 16408
rect 23615 16405 23627 16439
rect 23569 16399 23627 16405
rect 23750 16396 23756 16448
rect 23808 16436 23814 16448
rect 24673 16439 24731 16445
rect 24673 16436 24685 16439
rect 23808 16408 24685 16436
rect 23808 16396 23814 16408
rect 24673 16405 24685 16408
rect 24719 16405 24731 16439
rect 24673 16399 24731 16405
rect 25038 16396 25044 16448
rect 25096 16396 25102 16448
rect 25133 16439 25191 16445
rect 25133 16405 25145 16439
rect 25179 16436 25191 16439
rect 25314 16436 25320 16448
rect 25179 16408 25320 16436
rect 25179 16405 25191 16408
rect 25133 16399 25191 16405
rect 25314 16396 25320 16408
rect 25372 16396 25378 16448
rect 25406 16396 25412 16448
rect 25464 16436 25470 16448
rect 26620 16445 26648 16476
rect 25869 16439 25927 16445
rect 25869 16436 25881 16439
rect 25464 16408 25881 16436
rect 25464 16396 25470 16408
rect 25869 16405 25881 16408
rect 25915 16405 25927 16439
rect 25869 16399 25927 16405
rect 26605 16439 26663 16445
rect 26605 16405 26617 16439
rect 26651 16405 26663 16439
rect 26712 16436 26740 16544
rect 27706 16532 27712 16584
rect 27764 16572 27770 16584
rect 28169 16575 28227 16581
rect 28169 16572 28181 16575
rect 27764 16544 28181 16572
rect 27764 16532 27770 16544
rect 28169 16541 28181 16544
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 28261 16575 28319 16581
rect 28261 16541 28273 16575
rect 28307 16572 28319 16575
rect 28626 16572 28632 16584
rect 28307 16544 28632 16572
rect 28307 16541 28319 16544
rect 28261 16535 28319 16541
rect 28626 16532 28632 16544
rect 28684 16532 28690 16584
rect 26973 16507 27031 16513
rect 26973 16473 26985 16507
rect 27019 16504 27031 16507
rect 28442 16504 28448 16516
rect 27019 16476 28448 16504
rect 27019 16473 27031 16476
rect 26973 16467 27031 16473
rect 28442 16464 28448 16476
rect 28500 16464 28506 16516
rect 27801 16439 27859 16445
rect 27801 16436 27813 16439
rect 26712 16408 27813 16436
rect 26605 16399 26663 16405
rect 27801 16405 27813 16408
rect 27847 16405 27859 16439
rect 27801 16399 27859 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 4890 16192 4896 16244
rect 4948 16232 4954 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 4948 16204 7297 16232
rect 4948 16192 4954 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 7285 16195 7343 16201
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 10134 16232 10140 16244
rect 7432 16204 10140 16232
rect 7432 16192 7438 16204
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10226 16192 10232 16244
rect 10284 16192 10290 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 21450 16232 21456 16244
rect 12492 16204 21456 16232
rect 12492 16192 12498 16204
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 23753 16235 23811 16241
rect 23753 16201 23765 16235
rect 23799 16232 23811 16235
rect 24026 16232 24032 16244
rect 23799 16204 24032 16232
rect 23799 16201 23811 16204
rect 23753 16195 23811 16201
rect 24026 16192 24032 16204
rect 24084 16232 24090 16244
rect 24486 16232 24492 16244
rect 24084 16204 24492 16232
rect 24084 16192 24090 16204
rect 24486 16192 24492 16204
rect 24544 16192 24550 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 25004 16204 26617 16232
rect 25004 16192 25010 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 26786 16192 26792 16244
rect 26844 16232 26850 16244
rect 26973 16235 27031 16241
rect 26973 16232 26985 16235
rect 26844 16204 26985 16232
rect 26844 16192 26850 16204
rect 26973 16201 26985 16204
rect 27019 16201 27031 16235
rect 26973 16195 27031 16201
rect 27614 16192 27620 16244
rect 27672 16232 27678 16244
rect 27709 16235 27767 16241
rect 27709 16232 27721 16235
rect 27672 16204 27721 16232
rect 27672 16192 27678 16204
rect 27709 16201 27721 16204
rect 27755 16232 27767 16235
rect 28626 16232 28632 16244
rect 27755 16204 28632 16232
rect 27755 16201 27767 16204
rect 27709 16195 27767 16201
rect 28626 16192 28632 16204
rect 28684 16192 28690 16244
rect 3326 16124 3332 16176
rect 3384 16164 3390 16176
rect 4341 16167 4399 16173
rect 4341 16164 4353 16167
rect 3384 16136 4353 16164
rect 3384 16124 3390 16136
rect 4341 16133 4353 16136
rect 4387 16133 4399 16167
rect 4341 16127 4399 16133
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 8757 16167 8815 16173
rect 8757 16164 8769 16167
rect 5868 16136 8769 16164
rect 5868 16124 5874 16136
rect 8312 16108 8340 16136
rect 8757 16133 8769 16136
rect 8803 16133 8815 16167
rect 10594 16164 10600 16176
rect 9982 16136 10600 16164
rect 8757 16127 8815 16133
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 12250 16124 12256 16176
rect 12308 16124 12314 16176
rect 12710 16124 12716 16176
rect 12768 16124 12774 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 14568 16136 19717 16164
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1811 16068 2774 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2746 16028 2774 16068
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 3786 16056 3792 16108
rect 3844 16096 3850 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 3844 16068 5641 16096
rect 3844 16056 3850 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 7374 16096 7380 16108
rect 5629 16059 5687 16065
rect 5828 16068 7380 16096
rect 4062 16028 4068 16040
rect 2746 16000 4068 16028
rect 2041 15991 2099 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 5718 15988 5724 16040
rect 5776 15988 5782 16040
rect 5261 15963 5319 15969
rect 5261 15929 5273 15963
rect 5307 15960 5319 15963
rect 5828 15960 5856 16068
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 8294 16056 8300 16108
rect 8352 16056 8358 16108
rect 8478 16056 8484 16108
rect 8536 16056 8542 16108
rect 11146 16056 11152 16108
rect 11204 16056 11210 16108
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6178 16028 6184 16040
rect 5951 16000 6184 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6178 15988 6184 16000
rect 6236 16028 6242 16040
rect 6546 16028 6552 16040
rect 6236 16000 6552 16028
rect 6236 15988 6242 16000
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 6638 15988 6644 16040
rect 6696 15988 6702 16040
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7524 16000 7757 16028
rect 7524 15988 7530 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 7929 16031 7987 16037
rect 7929 15997 7941 16031
rect 7975 16028 7987 16031
rect 8202 16028 8208 16040
rect 7975 16000 8208 16028
rect 7975 15997 7987 16000
rect 7929 15991 7987 15997
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8312 16028 8340 16056
rect 9950 16028 9956 16040
rect 8312 16000 9956 16028
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 14568 16028 14596 16136
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 14642 16056 14648 16108
rect 14700 16056 14706 16108
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 16301 16099 16359 16105
rect 14792 16068 15608 16096
rect 14792 16056 14798 16068
rect 10468 16000 14596 16028
rect 14829 16031 14887 16037
rect 10468 15988 10474 16000
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 5307 15932 5856 15960
rect 9968 15960 9996 15988
rect 10318 15960 10324 15972
rect 9968 15932 10324 15960
rect 5307 15929 5319 15932
rect 5261 15923 5319 15929
rect 10318 15920 10324 15932
rect 10376 15960 10382 15972
rect 10870 15960 10876 15972
rect 10376 15932 10876 15960
rect 10376 15920 10382 15932
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 10962 15920 10968 15972
rect 11020 15920 11026 15972
rect 13630 15920 13636 15972
rect 13688 15960 13694 15972
rect 14844 15960 14872 15991
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 15160 16000 15485 16028
rect 15160 15988 15166 16000
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15580 16028 15608 16068
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 17586 16096 17592 16108
rect 16347 16068 17592 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 15580 16000 16804 16028
rect 15473 15991 15531 15997
rect 13688 15932 14872 15960
rect 13688 15920 13694 15932
rect 15286 15920 15292 15972
rect 15344 15960 15350 15972
rect 15930 15960 15936 15972
rect 15344 15932 15936 15960
rect 15344 15920 15350 15932
rect 15930 15920 15936 15932
rect 15988 15960 15994 15972
rect 16669 15963 16727 15969
rect 16669 15960 16681 15963
rect 15988 15932 16681 15960
rect 15988 15920 15994 15932
rect 16669 15929 16681 15932
rect 16715 15929 16727 15963
rect 16669 15923 16727 15929
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 8570 15892 8576 15904
rect 5684 15864 8576 15892
rect 5684 15852 5690 15864
rect 8570 15852 8576 15864
rect 8628 15892 8634 15904
rect 12066 15892 12072 15904
rect 8628 15864 12072 15892
rect 8628 15852 8634 15864
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12894 15852 12900 15904
rect 12952 15892 12958 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 12952 15864 13737 15892
rect 12952 15852 12958 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 13725 15855 13783 15861
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13964 15864 14289 15892
rect 13964 15852 13970 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 16114 15852 16120 15904
rect 16172 15852 16178 15904
rect 16776 15892 16804 16000
rect 16850 15988 16856 16040
rect 16908 16028 16914 16040
rect 17788 16028 17816 16059
rect 17862 16056 17868 16108
rect 17920 16056 17926 16108
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 19150 16096 19156 16108
rect 18647 16068 19156 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19720 16096 19748 16127
rect 20438 16124 20444 16176
rect 20496 16124 20502 16176
rect 21818 16164 21824 16176
rect 20732 16136 21824 16164
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 19720 16068 20545 16096
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 16908 16000 17816 16028
rect 17880 16000 17969 16028
rect 16908 15988 16914 16000
rect 17310 15920 17316 15972
rect 17368 15960 17374 15972
rect 17405 15963 17463 15969
rect 17405 15960 17417 15963
rect 17368 15932 17417 15960
rect 17368 15920 17374 15932
rect 17405 15929 17417 15932
rect 17451 15929 17463 15963
rect 17405 15923 17463 15929
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 17880 15960 17908 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 18874 15988 18880 16040
rect 18932 15988 18938 16040
rect 20732 16037 20760 16136
rect 21818 16124 21824 16136
rect 21876 16124 21882 16176
rect 23474 16124 23480 16176
rect 23532 16164 23538 16176
rect 23661 16167 23719 16173
rect 23661 16164 23673 16167
rect 23532 16136 23673 16164
rect 23532 16124 23538 16136
rect 23661 16133 23673 16136
rect 23707 16164 23719 16167
rect 24394 16164 24400 16176
rect 23707 16136 24400 16164
rect 23707 16133 23719 16136
rect 23661 16127 23719 16133
rect 24394 16124 24400 16136
rect 24452 16124 24458 16176
rect 25038 16124 25044 16176
rect 25096 16164 25102 16176
rect 25406 16164 25412 16176
rect 25096 16136 25412 16164
rect 25096 16124 25102 16136
rect 25406 16124 25412 16136
rect 25464 16124 25470 16176
rect 26804 16164 26832 16192
rect 26358 16136 26832 16164
rect 22281 16099 22339 16105
rect 21453 16083 21511 16089
rect 21453 16049 21465 16083
rect 21499 16049 21511 16083
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22922 16096 22928 16108
rect 22327 16068 22928 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 21453 16043 21511 16049
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 17552 15932 17908 15960
rect 20073 15963 20131 15969
rect 17552 15920 17558 15932
rect 20073 15929 20085 15963
rect 20119 15960 20131 15963
rect 21358 15960 21364 15972
rect 20119 15932 21364 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 21468 15960 21496 16043
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21784 16000 22017 16028
rect 21784 15988 21790 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 23937 16031 23995 16037
rect 23937 15997 23949 16031
rect 23983 16028 23995 16031
rect 24026 16028 24032 16040
rect 23983 16000 24032 16028
rect 23983 15997 23995 16000
rect 23937 15991 23995 15997
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 25130 15988 25136 16040
rect 25188 16028 25194 16040
rect 27246 16028 27252 16040
rect 25188 16000 27252 16028
rect 25188 15988 25194 16000
rect 27246 15988 27252 16000
rect 27304 15988 27310 16040
rect 21468 15932 23796 15960
rect 16942 15892 16948 15904
rect 16776 15864 16948 15892
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 18598 15892 18604 15904
rect 17184 15864 18604 15892
rect 17184 15852 17190 15864
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 20806 15892 20812 15904
rect 19668 15864 20812 15892
rect 19668 15852 19674 15864
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 21542 15852 21548 15904
rect 21600 15892 21606 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 21600 15864 23305 15892
rect 21600 15852 21606 15864
rect 23293 15861 23305 15864
rect 23339 15861 23351 15895
rect 23768 15892 23796 15932
rect 23842 15920 23848 15972
rect 23900 15960 23906 15972
rect 29730 15960 29736 15972
rect 23900 15932 24624 15960
rect 23900 15920 23906 15932
rect 24302 15892 24308 15904
rect 23768 15864 24308 15892
rect 23293 15855 23351 15861
rect 24302 15852 24308 15864
rect 24360 15852 24366 15904
rect 24596 15892 24624 15932
rect 26160 15932 29736 15960
rect 26160 15892 26188 15932
rect 29730 15920 29736 15932
rect 29788 15920 29794 15972
rect 24596 15864 26188 15892
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7248 15660 7849 15688
rect 7248 15648 7254 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8720 15660 9321 15688
rect 8720 15648 8726 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 12802 15688 12808 15700
rect 11020 15660 12808 15688
rect 11020 15648 11026 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13173 15691 13231 15697
rect 13173 15657 13185 15691
rect 13219 15688 13231 15691
rect 13354 15688 13360 15700
rect 13219 15660 13360 15688
rect 13219 15657 13231 15660
rect 13173 15651 13231 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 23934 15688 23940 15700
rect 13740 15660 23940 15688
rect 6178 15620 6184 15632
rect 4632 15592 6184 15620
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 4632 15561 4660 15592
rect 6178 15580 6184 15592
rect 6236 15580 6242 15632
rect 7558 15620 7564 15632
rect 7300 15592 7564 15620
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5592 15524 5641 15552
rect 5592 15512 5598 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3418 15484 3424 15496
rect 1811 15456 3424 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 5828 15484 5856 15515
rect 6822 15512 6828 15564
rect 6880 15512 6886 15564
rect 6914 15512 6920 15564
rect 6972 15512 6978 15564
rect 7190 15484 7196 15496
rect 5828 15456 7196 15484
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 5537 15419 5595 15425
rect 5537 15416 5549 15419
rect 3988 15388 5549 15416
rect 3988 15357 4016 15388
rect 5537 15385 5549 15388
rect 5583 15385 5595 15419
rect 5537 15379 5595 15385
rect 6733 15419 6791 15425
rect 6733 15385 6745 15419
rect 6779 15416 6791 15419
rect 7300 15416 7328 15592
rect 7558 15580 7564 15592
rect 7616 15580 7622 15632
rect 9646 15592 10088 15620
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 8352 15524 8401 15552
rect 8352 15512 8358 15524
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 9214 15512 9220 15564
rect 9272 15552 9278 15564
rect 9646 15552 9674 15592
rect 9272 15524 9674 15552
rect 10060 15552 10088 15592
rect 10336 15592 11560 15620
rect 10336 15552 10364 15592
rect 10060 15524 10364 15552
rect 9272 15512 9278 15524
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 10928 15524 11437 15552
rect 10928 15512 10934 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11532 15552 11560 15592
rect 12066 15580 12072 15632
rect 12124 15580 12130 15632
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 13541 15623 13599 15629
rect 13541 15620 13553 15623
rect 12216 15592 13553 15620
rect 12216 15580 12222 15592
rect 13541 15589 13553 15592
rect 13587 15589 13599 15623
rect 13541 15583 13599 15589
rect 12713 15555 12771 15561
rect 11532 15524 12572 15552
rect 11425 15515 11483 15521
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 12437 15487 12495 15493
rect 12437 15484 12449 15487
rect 8720 15456 12449 15484
rect 8720 15444 8726 15456
rect 12437 15453 12449 15456
rect 12483 15453 12495 15487
rect 12544 15484 12572 15524
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12894 15552 12900 15564
rect 12759 15524 12900 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13630 15484 13636 15496
rect 12544 15456 13636 15484
rect 12437 15447 12495 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 13740 15493 13768 15660
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 24486 15648 24492 15700
rect 24544 15648 24550 15700
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 14461 15623 14519 15629
rect 14461 15620 14473 15623
rect 13872 15592 14473 15620
rect 13872 15580 13878 15592
rect 14461 15589 14473 15592
rect 14507 15589 14519 15623
rect 14461 15583 14519 15589
rect 15838 15580 15844 15632
rect 15896 15580 15902 15632
rect 21726 15620 21732 15632
rect 21652 15592 21732 15620
rect 15010 15512 15016 15564
rect 15068 15512 15074 15564
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 15102 15484 15108 15496
rect 14875 15456 15108 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 6779 15388 7328 15416
rect 6779 15385 6791 15388
rect 6733 15379 6791 15385
rect 7558 15376 7564 15428
rect 7616 15416 7622 15428
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 7616 15388 8309 15416
rect 7616 15376 7622 15388
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9769 15419 9827 15425
rect 9769 15416 9781 15419
rect 9272 15388 9781 15416
rect 9272 15376 9278 15388
rect 9769 15385 9781 15388
rect 9815 15416 9827 15419
rect 9858 15416 9864 15428
rect 9815 15388 9864 15416
rect 9815 15385 9827 15388
rect 9769 15379 9827 15385
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 9950 15376 9956 15428
rect 10008 15376 10014 15428
rect 10229 15419 10287 15425
rect 10229 15385 10241 15419
rect 10275 15416 10287 15419
rect 10962 15416 10968 15428
rect 10275 15388 10968 15416
rect 10275 15385 10287 15388
rect 10229 15379 10287 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11241 15419 11299 15425
rect 11241 15416 11253 15419
rect 11112 15388 11253 15416
rect 11112 15376 11118 15388
rect 11241 15385 11253 15388
rect 11287 15416 11299 15419
rect 11287 15388 12664 15416
rect 11287 15385 11299 15388
rect 11241 15379 11299 15385
rect 3973 15351 4031 15357
rect 3973 15317 3985 15351
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 4338 15308 4344 15360
rect 4396 15308 4402 15360
rect 4433 15351 4491 15357
rect 4433 15317 4445 15351
rect 4479 15348 4491 15351
rect 4798 15348 4804 15360
rect 4479 15320 4804 15348
rect 4479 15317 4491 15320
rect 4433 15311 4491 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 6362 15308 6368 15360
rect 6420 15308 6426 15360
rect 7466 15308 7472 15360
rect 7524 15308 7530 15360
rect 7834 15308 7840 15360
rect 7892 15348 7898 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7892 15320 8217 15348
rect 7892 15308 7898 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8205 15311 8263 15317
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 10410 15348 10416 15360
rect 8720 15320 10416 15348
rect 8720 15308 8726 15320
rect 10410 15308 10416 15320
rect 10468 15308 10474 15360
rect 10870 15308 10876 15360
rect 10928 15308 10934 15360
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11790 15348 11796 15360
rect 11379 15320 11796 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 12636 15348 12664 15388
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 15473 15419 15531 15425
rect 15473 15416 15485 15419
rect 13320 15388 15485 15416
rect 13320 15376 13326 15388
rect 15473 15385 15485 15388
rect 15519 15416 15531 15419
rect 16209 15419 16267 15425
rect 16209 15416 16221 15419
rect 15519 15388 16221 15416
rect 15519 15385 15531 15388
rect 15473 15379 15531 15385
rect 16209 15385 16221 15388
rect 16255 15385 16267 15419
rect 16500 15416 16528 15515
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19484 15524 20269 15552
rect 19484 15512 19490 15524
rect 20257 15521 20269 15524
rect 20303 15552 20315 15555
rect 20622 15552 20628 15564
rect 20303 15524 20628 15552
rect 20303 15521 20315 15524
rect 20257 15515 20315 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 19610 15444 19616 15496
rect 19668 15444 19674 15496
rect 21652 15470 21680 15592
rect 21726 15580 21732 15592
rect 21784 15620 21790 15632
rect 21910 15620 21916 15632
rect 21784 15592 21916 15620
rect 21784 15580 21790 15592
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 22094 15580 22100 15632
rect 22152 15620 22158 15632
rect 22741 15623 22799 15629
rect 22741 15620 22753 15623
rect 22152 15592 22753 15620
rect 22152 15580 22158 15592
rect 22741 15589 22753 15592
rect 22787 15589 22799 15623
rect 22741 15583 22799 15589
rect 21836 15524 22692 15552
rect 17310 15416 17316 15428
rect 16500 15388 17316 15416
rect 16209 15379 16267 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17770 15376 17776 15428
rect 17828 15376 17834 15428
rect 18598 15376 18604 15428
rect 18656 15416 18662 15428
rect 18656 15388 19472 15416
rect 18656 15376 18662 15388
rect 13354 15348 13360 15360
rect 12636 15320 13360 15348
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 14550 15308 14556 15360
rect 14608 15348 14614 15360
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 14608 15320 14933 15348
rect 14608 15308 14614 15320
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 14921 15311 14979 15317
rect 15378 15308 15384 15360
rect 15436 15348 15442 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 15436 15320 16313 15348
rect 15436 15308 15442 15320
rect 16301 15317 16313 15320
rect 16347 15348 16359 15351
rect 16574 15348 16580 15360
rect 16347 15320 16580 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 19444 15357 19472 15388
rect 19886 15376 19892 15428
rect 19944 15416 19950 15428
rect 20533 15419 20591 15425
rect 20533 15416 20545 15419
rect 19944 15388 20545 15416
rect 19944 15376 19950 15388
rect 20533 15385 20545 15388
rect 20579 15385 20591 15419
rect 20533 15379 20591 15385
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 17460 15320 18797 15348
rect 17460 15308 17466 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 19429 15351 19487 15357
rect 19429 15317 19441 15351
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 19702 15308 19708 15360
rect 19760 15348 19766 15360
rect 20438 15348 20444 15360
rect 19760 15320 20444 15348
rect 19760 15308 19766 15320
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 20548 15348 20576 15379
rect 21836 15348 21864 15524
rect 21910 15444 21916 15496
rect 21968 15484 21974 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 21968 15456 22293 15484
rect 21968 15444 21974 15456
rect 22281 15453 22293 15456
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 20548 15320 21864 15348
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21968 15320 22017 15348
rect 21968 15308 21974 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22296 15348 22324 15447
rect 22664 15416 22692 15524
rect 22756 15484 22784 15583
rect 24302 15512 24308 15564
rect 24360 15552 24366 15564
rect 25222 15552 25228 15564
rect 24360 15524 25228 15552
rect 24360 15512 24366 15524
rect 25222 15512 25228 15524
rect 25280 15552 25286 15564
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 25280 15524 25789 15552
rect 25280 15512 25286 15524
rect 25777 15521 25789 15524
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22756 15456 23121 15484
rect 23109 15453 23121 15456
rect 23155 15484 23167 15487
rect 23290 15484 23296 15496
rect 23155 15456 23296 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 26050 15444 26056 15496
rect 26108 15484 26114 15496
rect 26108 15456 31754 15484
rect 26108 15444 26114 15456
rect 23566 15416 23572 15428
rect 22664 15388 23572 15416
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 23934 15376 23940 15428
rect 23992 15376 23998 15428
rect 26142 15416 26148 15428
rect 25608 15388 26148 15416
rect 25608 15360 25636 15388
rect 26142 15376 26148 15388
rect 26200 15416 26206 15428
rect 26237 15419 26295 15425
rect 26237 15416 26249 15419
rect 26200 15388 26249 15416
rect 26200 15376 26206 15388
rect 26237 15385 26249 15388
rect 26283 15416 26295 15419
rect 31726 15416 31754 15456
rect 48682 15416 48688 15428
rect 26283 15388 29040 15416
rect 31726 15388 48688 15416
rect 26283 15385 26295 15388
rect 26237 15379 26295 15385
rect 22738 15348 22744 15360
rect 22296 15320 22744 15348
rect 22005 15311 22063 15317
rect 22738 15308 22744 15320
rect 22796 15348 22802 15360
rect 23842 15348 23848 15360
rect 22796 15320 23848 15348
rect 22796 15308 22802 15320
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 25222 15308 25228 15360
rect 25280 15308 25286 15360
rect 25590 15308 25596 15360
rect 25648 15308 25654 15360
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15348 25743 15351
rect 26050 15348 26056 15360
rect 25731 15320 26056 15348
rect 25731 15317 25743 15320
rect 25685 15311 25743 15317
rect 26050 15308 26056 15320
rect 26108 15348 26114 15360
rect 26421 15351 26479 15357
rect 26421 15348 26433 15351
rect 26108 15320 26433 15348
rect 26108 15308 26114 15320
rect 26421 15317 26433 15320
rect 26467 15317 26479 15351
rect 29012 15348 29040 15388
rect 48682 15376 48688 15388
rect 48740 15376 48746 15428
rect 49234 15348 49240 15360
rect 29012 15320 49240 15348
rect 26421 15311 26479 15317
rect 49234 15308 49240 15320
rect 49292 15308 49298 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 4120 15116 6745 15144
rect 4120 15104 4126 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 8662 15144 8668 15156
rect 6972 15116 8668 15144
rect 6972 15104 6978 15116
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 11238 15144 11244 15156
rect 9631 15116 11244 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12676 15116 13001 15144
rect 12676 15104 12682 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 16666 15144 16672 15156
rect 13136 15116 16672 15144
rect 13136 15104 13142 15116
rect 16666 15104 16672 15116
rect 16724 15104 16730 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 22094 15144 22100 15156
rect 18472 15116 22100 15144
rect 18472 15104 18478 15116
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 23566 15104 23572 15156
rect 23624 15144 23630 15156
rect 23753 15147 23811 15153
rect 23753 15144 23765 15147
rect 23624 15116 23765 15144
rect 23624 15104 23630 15116
rect 23753 15113 23765 15116
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 23842 15104 23848 15156
rect 23900 15144 23906 15156
rect 24029 15147 24087 15153
rect 24029 15144 24041 15147
rect 23900 15116 24041 15144
rect 23900 15104 23906 15116
rect 24029 15113 24041 15116
rect 24075 15144 24087 15147
rect 24213 15147 24271 15153
rect 24213 15144 24225 15147
rect 24075 15116 24225 15144
rect 24075 15113 24087 15116
rect 24029 15107 24087 15113
rect 24213 15113 24225 15116
rect 24259 15113 24271 15147
rect 24213 15107 24271 15113
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 26786 15104 26792 15156
rect 26844 15144 26850 15156
rect 26973 15147 27031 15153
rect 26973 15144 26985 15147
rect 26844 15116 26985 15144
rect 26844 15104 26850 15116
rect 26973 15113 26985 15116
rect 27019 15113 27031 15147
rect 26973 15107 27031 15113
rect 4433 15079 4491 15085
rect 1780 15048 4108 15076
rect 1780 15017 1808 15048
rect 4080 15020 4108 15048
rect 4433 15045 4445 15079
rect 4479 15076 4491 15079
rect 4706 15076 4712 15088
rect 4479 15048 4712 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 6270 15076 6276 15088
rect 5658 15048 6276 15076
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 7653 15079 7711 15085
rect 7653 15045 7665 15079
rect 7699 15076 7711 15079
rect 7742 15076 7748 15088
rect 7699 15048 7748 15076
rect 7699 15045 7711 15048
rect 7653 15039 7711 15045
rect 7742 15036 7748 15048
rect 7800 15036 7806 15088
rect 8570 15036 8576 15088
rect 8628 15036 8634 15088
rect 8757 15079 8815 15085
rect 8757 15045 8769 15079
rect 8803 15076 8815 15079
rect 8846 15076 8852 15088
rect 8803 15048 8852 15076
rect 8803 15045 8815 15048
rect 8757 15039 8815 15045
rect 8846 15036 8852 15048
rect 8904 15036 8910 15088
rect 9030 15036 9036 15088
rect 9088 15076 9094 15088
rect 9677 15079 9735 15085
rect 9677 15076 9689 15079
rect 9088 15048 9689 15076
rect 9088 15036 9094 15048
rect 9677 15045 9689 15048
rect 9723 15045 9735 15079
rect 9677 15039 9735 15045
rect 9858 15036 9864 15088
rect 9916 15036 9922 15088
rect 10778 15036 10784 15088
rect 10836 15036 10842 15088
rect 13262 15076 13268 15088
rect 10888 15048 13268 15076
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 3712 14940 3740 14971
rect 4062 14968 4068 15020
rect 4120 14968 4126 15020
rect 4154 14968 4160 15020
rect 4212 14968 4218 15020
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 6178 15008 6184 15020
rect 5868 14980 6184 15008
rect 5868 14968 5874 14980
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 15008 6699 15011
rect 7392 15008 7512 15012
rect 9876 15008 9904 15036
rect 6687 14984 9904 15008
rect 6687 14980 7420 14984
rect 7484 14980 9904 14984
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10888 15017 10916 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 13449 15079 13507 15085
rect 13449 15045 13461 15079
rect 13495 15076 13507 15079
rect 14093 15079 14151 15085
rect 14093 15076 14105 15079
rect 13495 15048 14105 15076
rect 13495 15045 13507 15048
rect 13449 15039 13507 15045
rect 14093 15045 14105 15048
rect 14139 15076 14151 15079
rect 14734 15076 14740 15088
rect 14139 15048 14740 15076
rect 14139 15045 14151 15048
rect 14093 15039 14151 15045
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 14829 15079 14887 15085
rect 14829 15045 14841 15079
rect 14875 15076 14887 15079
rect 15102 15076 15108 15088
rect 14875 15048 15108 15076
rect 14875 15045 14887 15048
rect 14829 15039 14887 15045
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 15286 15036 15292 15088
rect 15344 15036 15350 15088
rect 16574 15036 16580 15088
rect 16632 15076 16638 15088
rect 16761 15079 16819 15085
rect 16761 15076 16773 15079
rect 16632 15048 16773 15076
rect 16632 15036 16638 15048
rect 16761 15045 16773 15048
rect 16807 15076 16819 15079
rect 19518 15076 19524 15088
rect 16807 15048 19524 15076
rect 16807 15045 16819 15048
rect 16761 15039 16819 15045
rect 19518 15036 19524 15048
rect 19576 15036 19582 15088
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 21634 15076 21640 15088
rect 20211 15048 21640 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 22738 15036 22744 15088
rect 22796 15036 22802 15088
rect 24964 15076 24992 15104
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 24964 15048 25145 15076
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 26804 15076 26832 15104
rect 26358 15048 26832 15076
rect 25133 15039 25191 15045
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 10008 14980 10885 15008
rect 10008 14968 10014 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 12124 14980 13369 15008
rect 12124 14968 12130 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 17586 14968 17592 15020
rect 17644 15008 17650 15020
rect 19702 15008 19708 15020
rect 17644 14980 19708 15008
rect 17644 14968 17650 14980
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 20036 14980 20085 15008
rect 20036 14968 20042 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20180 14980 20484 15008
rect 7282 14940 7288 14952
rect 3712 14912 7288 14940
rect 2041 14903 2099 14909
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 7650 14900 7656 14952
rect 7708 14940 7714 14952
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 7708 14912 7757 14940
rect 7708 14900 7714 14912
rect 7745 14909 7757 14912
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 3602 14832 3608 14884
rect 3660 14872 3666 14884
rect 4062 14872 4068 14884
rect 3660 14844 4068 14872
rect 3660 14832 3666 14844
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 4488 14776 5917 14804
rect 4488 14764 4494 14776
rect 5905 14773 5917 14776
rect 5951 14804 5963 14807
rect 6822 14804 6828 14816
rect 5951 14776 6828 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 7760 14804 7788 14903
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 9858 14900 9864 14952
rect 9916 14900 9922 14952
rect 10965 14943 11023 14949
rect 10152 14912 10364 14940
rect 8294 14832 8300 14884
rect 8352 14872 8358 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 8352 14844 9229 14872
rect 8352 14832 8358 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 10152 14872 10180 14912
rect 9548 14844 10180 14872
rect 10336 14872 10364 14912
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11330 14940 11336 14952
rect 11011 14912 11336 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 12250 14900 12256 14952
rect 12308 14940 12314 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 12308 14912 13553 14940
rect 12308 14900 12314 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13556 14872 13584 14903
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 14332 14912 14565 14940
rect 14332 14900 14338 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 16114 14940 16120 14952
rect 14553 14903 14611 14909
rect 14660 14912 16120 14940
rect 13722 14872 13728 14884
rect 10336 14844 10826 14872
rect 13556 14844 13728 14872
rect 9548 14832 9554 14844
rect 10042 14804 10048 14816
rect 7760 14776 10048 14804
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 10798 14804 10826 14844
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 14660 14872 14688 14912
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 20180 14940 20208 14980
rect 19300 14912 19840 14940
rect 19300 14900 19306 14912
rect 13832 14844 14688 14872
rect 13832 14804 13860 14844
rect 15838 14832 15844 14884
rect 15896 14872 15902 14884
rect 17586 14872 17592 14884
rect 15896 14844 17592 14872
rect 15896 14832 15902 14844
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 19610 14872 19616 14884
rect 17920 14844 19616 14872
rect 17920 14832 17926 14844
rect 19610 14832 19616 14844
rect 19668 14832 19674 14884
rect 19702 14832 19708 14884
rect 19760 14832 19766 14884
rect 19812 14872 19840 14912
rect 19996 14912 20208 14940
rect 20349 14943 20407 14949
rect 19996 14872 20024 14912
rect 20349 14909 20361 14943
rect 20395 14909 20407 14943
rect 20456 14940 20484 14980
rect 20622 14968 20628 15020
rect 20680 15008 20686 15020
rect 22002 15008 22008 15020
rect 20680 14980 22008 15008
rect 20680 14968 20686 14980
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 23992 14980 24869 15008
rect 23992 14968 23998 14980
rect 24857 14977 24869 14980
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20456 14912 20913 14940
rect 20349 14903 20407 14909
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14940 22339 14943
rect 22646 14940 22652 14952
rect 22327 14912 22652 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 19812 14844 20024 14872
rect 20364 14872 20392 14903
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 21910 14872 21916 14884
rect 20364 14844 21916 14872
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 24854 14872 24860 14884
rect 23768 14844 24860 14872
rect 10798 14776 13860 14804
rect 14182 14764 14188 14816
rect 14240 14804 14246 14816
rect 15286 14804 15292 14816
rect 14240 14776 15292 14804
rect 14240 14764 14246 14776
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 16298 14764 16304 14816
rect 16356 14764 16362 14816
rect 17770 14764 17776 14816
rect 17828 14804 17834 14816
rect 18874 14804 18880 14816
rect 17828 14776 18880 14804
rect 17828 14764 17834 14776
rect 18874 14764 18880 14776
rect 18932 14804 18938 14816
rect 19153 14807 19211 14813
rect 19153 14804 19165 14807
rect 18932 14776 19165 14804
rect 18932 14764 18938 14776
rect 19153 14773 19165 14776
rect 19199 14773 19211 14807
rect 19153 14767 19211 14773
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 23768 14804 23796 14844
rect 24854 14832 24860 14844
rect 24912 14832 24918 14884
rect 19576 14776 23796 14804
rect 19576 14764 19582 14776
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4212 14572 4261 14600
rect 4212 14560 4218 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 4890 14600 4896 14612
rect 4764 14572 4896 14600
rect 4764 14560 4770 14572
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 9214 14600 9220 14612
rect 5040 14572 9220 14600
rect 5040 14560 5046 14572
rect 9214 14560 9220 14572
rect 9272 14560 9278 14612
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 10686 14600 10692 14612
rect 9447 14572 10692 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 10836 14572 11621 14600
rect 10836 14560 10842 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 13538 14600 13544 14612
rect 11609 14563 11667 14569
rect 11716 14572 13544 14600
rect 7190 14492 7196 14544
rect 7248 14532 7254 14544
rect 7650 14532 7656 14544
rect 7248 14504 7656 14532
rect 7248 14492 7254 14504
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 9858 14532 9864 14544
rect 8496 14504 9864 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 4246 14424 4252 14476
rect 4304 14424 4310 14476
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 4488 14436 4813 14464
rect 4488 14424 4494 14436
rect 4801 14433 4813 14436
rect 4847 14433 4859 14467
rect 4801 14427 4859 14433
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 8496 14473 8524 14504
rect 9858 14492 9864 14504
rect 9916 14532 9922 14544
rect 10042 14532 10048 14544
rect 9916 14504 10048 14532
rect 9916 14492 9922 14504
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 10192 14504 10364 14532
rect 10192 14492 10198 14504
rect 8481 14467 8539 14473
rect 6788 14436 8248 14464
rect 6788 14424 6794 14436
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 4264 14396 4292 14424
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 1811 14368 2774 14396
rect 4264 14368 4629 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 2746 14328 2774 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5224 14368 5457 14396
rect 5224 14356 5230 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7834 14396 7840 14408
rect 7248 14368 7840 14396
rect 7248 14356 7254 14368
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 8220 14405 8248 14436
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 9674 14464 9680 14476
rect 8720 14436 9680 14464
rect 8720 14424 8726 14436
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9953 14467 10011 14473
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10226 14464 10232 14476
rect 9999 14436 10232 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10336 14464 10364 14504
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10336 14436 11161 14464
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 9766 14396 9772 14408
rect 8343 14368 9772 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10870 14396 10876 14408
rect 9907 14368 10876 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 5721 14331 5779 14337
rect 2746 14300 4844 14328
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 4212 14232 4721 14260
rect 4212 14220 4218 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 4816 14260 4844 14300
rect 5721 14297 5733 14331
rect 5767 14328 5779 14331
rect 5810 14328 5816 14340
rect 5767 14300 5816 14328
rect 5767 14297 5779 14300
rect 5721 14291 5779 14297
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 6270 14288 6276 14340
rect 6328 14288 6334 14340
rect 9398 14328 9404 14340
rect 7024 14300 9404 14328
rect 7024 14260 7052 14300
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 10134 14328 10140 14340
rect 9732 14300 10140 14328
rect 9732 14288 9738 14300
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10226 14288 10232 14340
rect 10284 14328 10290 14340
rect 11716 14328 11744 14572
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13722 14560 13728 14612
rect 13780 14560 13786 14612
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 14458 14600 14464 14612
rect 14415 14572 14464 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 15102 14560 15108 14612
rect 15160 14600 15166 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 15160 14572 18613 14600
rect 15160 14560 15166 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 18874 14560 18880 14612
rect 18932 14560 18938 14612
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 21729 14603 21787 14609
rect 21729 14600 21741 14603
rect 21140 14572 21741 14600
rect 21140 14560 21146 14572
rect 21729 14569 21741 14572
rect 21775 14569 21787 14603
rect 34882 14600 34888 14612
rect 21729 14563 21787 14569
rect 22066 14572 34888 14600
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14532 19487 14535
rect 22066 14532 22094 14572
rect 34882 14560 34888 14572
rect 34940 14560 34946 14612
rect 19475 14504 22094 14532
rect 19475 14501 19487 14504
rect 19429 14495 19487 14501
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12802 14464 12808 14476
rect 12308 14436 12808 14464
rect 12308 14424 12314 14436
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 12894 14424 12900 14476
rect 12952 14464 12958 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 12952 14436 14105 14464
rect 12952 14424 12958 14436
rect 14093 14433 14105 14436
rect 14139 14464 14151 14467
rect 14182 14464 14188 14476
rect 14139 14436 14188 14464
rect 14139 14433 14151 14436
rect 14093 14427 14151 14433
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 16298 14464 16304 14476
rect 14967 14436 16304 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14464 16911 14467
rect 17126 14464 17132 14476
rect 16899 14436 17132 14464
rect 16899 14433 16911 14436
rect 16853 14427 16911 14433
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 18322 14464 18328 14476
rect 17276 14436 18328 14464
rect 17276 14424 17282 14436
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 19300 14436 21097 14464
rect 19300 14424 19306 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22060 14436 22293 14464
rect 22060 14424 22066 14436
rect 22281 14433 22293 14436
rect 22327 14464 22339 14467
rect 23934 14464 23940 14476
rect 22327 14436 23940 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14464 25191 14467
rect 26329 14467 26387 14473
rect 26329 14464 26341 14467
rect 25179 14436 26341 14464
rect 25179 14433 25191 14436
rect 25133 14427 25191 14433
rect 26329 14433 26341 14436
rect 26375 14464 26387 14467
rect 26602 14464 26608 14476
rect 26375 14436 26608 14464
rect 26375 14433 26387 14436
rect 26329 14427 26387 14433
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 14332 14368 14657 14396
rect 14332 14356 14338 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 14645 14359 14703 14365
rect 18432 14368 19625 14396
rect 10284 14300 11744 14328
rect 10284 14288 10290 14300
rect 4816 14232 7052 14260
rect 4709 14223 4767 14229
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8812 14232 8953 14260
rect 8812 14220 8818 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9766 14220 9772 14272
rect 9824 14220 9830 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 11072 14269 11100 14300
rect 12250 14288 12256 14340
rect 12308 14288 12314 14340
rect 12710 14288 12716 14340
rect 12768 14288 12774 14340
rect 13556 14300 14412 14328
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 9916 14232 10609 14260
rect 9916 14220 9922 14232
rect 10597 14229 10609 14232
rect 10643 14229 10655 14263
rect 10597 14223 10655 14229
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13556 14260 13584 14300
rect 13228 14232 13584 14260
rect 14384 14260 14412 14300
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 16850 14328 16856 14340
rect 16224 14300 16856 14328
rect 16224 14260 16252 14300
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17129 14331 17187 14337
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17402 14328 17408 14340
rect 17175 14300 17408 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 17862 14288 17868 14340
rect 17920 14288 17926 14340
rect 14384 14232 16252 14260
rect 13228 14220 13234 14232
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 18432 14260 18460 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 25148 14396 25176 14427
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 19613 14359 19671 14365
rect 23952 14368 25176 14396
rect 20993 14331 21051 14337
rect 20993 14297 21005 14331
rect 21039 14328 21051 14331
rect 21082 14328 21088 14340
rect 21039 14300 21088 14328
rect 21039 14297 21051 14300
rect 20993 14291 21051 14297
rect 21082 14288 21088 14300
rect 21140 14288 21146 14340
rect 21910 14288 21916 14340
rect 21968 14328 21974 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 21968 14300 22569 14328
rect 21968 14288 21974 14300
rect 22557 14297 22569 14300
rect 22603 14297 22615 14331
rect 23842 14328 23848 14340
rect 23782 14300 23848 14328
rect 22557 14291 22615 14297
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 16540 14232 18460 14260
rect 16540 14220 16546 14232
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 21450 14260 21456 14272
rect 20947 14232 21456 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 21450 14220 21456 14232
rect 21508 14260 21514 14272
rect 21637 14263 21695 14269
rect 21637 14260 21649 14263
rect 21508 14232 21649 14260
rect 21508 14220 21514 14232
rect 21637 14229 21649 14232
rect 21683 14260 21695 14263
rect 21818 14260 21824 14272
rect 21683 14232 21824 14260
rect 21683 14229 21695 14232
rect 21637 14223 21695 14229
rect 21818 14220 21824 14232
rect 21876 14220 21882 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 23952 14260 23980 14368
rect 26142 14356 26148 14408
rect 26200 14396 26206 14408
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26200 14368 26985 14396
rect 26200 14356 26206 14368
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 24946 14288 24952 14340
rect 25004 14288 25010 14340
rect 25038 14288 25044 14340
rect 25096 14328 25102 14340
rect 25314 14328 25320 14340
rect 25096 14300 25320 14328
rect 25096 14288 25102 14300
rect 25314 14288 25320 14300
rect 25372 14288 25378 14340
rect 22796 14232 23980 14260
rect 24029 14263 24087 14269
rect 22796 14220 22802 14232
rect 24029 14229 24041 14263
rect 24075 14260 24087 14263
rect 24302 14260 24308 14272
rect 24075 14232 24308 14260
rect 24075 14229 24087 14232
rect 24029 14223 24087 14229
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 24964 14260 24992 14288
rect 25682 14260 25688 14272
rect 24964 14232 25688 14260
rect 25682 14220 25688 14232
rect 25740 14220 25746 14272
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 26142 14220 26148 14272
rect 26200 14260 26206 14272
rect 26237 14263 26295 14269
rect 26237 14260 26249 14263
rect 26200 14232 26249 14260
rect 26200 14220 26206 14232
rect 26237 14229 26249 14232
rect 26283 14260 26295 14263
rect 26789 14263 26847 14269
rect 26789 14260 26801 14263
rect 26283 14232 26801 14260
rect 26283 14229 26295 14232
rect 26237 14223 26295 14229
rect 26789 14229 26801 14232
rect 26835 14229 26847 14263
rect 26789 14223 26847 14229
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4154 14056 4160 14068
rect 4111 14028 4160 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 4982 14056 4988 14068
rect 4479 14028 4988 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6362 14056 6368 14068
rect 5675 14028 6368 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 4246 13948 4252 14000
rect 4304 13988 4310 14000
rect 5721 13991 5779 13997
rect 5721 13988 5733 13991
rect 4304 13960 5733 13988
rect 4304 13948 4310 13960
rect 5721 13957 5733 13960
rect 5767 13957 5779 13991
rect 6932 13988 6960 14019
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 7374 14016 7380 14068
rect 7432 14016 7438 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 9214 14056 9220 14068
rect 8159 14028 9220 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11480 14028 11621 14056
rect 11480 14016 11486 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 11609 14019 11667 14025
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 6932 13960 8493 13988
rect 5721 13951 5779 13957
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 10594 13948 10600 14000
rect 10652 13948 10658 14000
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 5626 13920 5632 13932
rect 3651 13892 5632 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 6328 13892 6377 13920
rect 6328 13880 6334 13892
rect 6365 13889 6377 13892
rect 6411 13920 6423 13923
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6411 13892 6561 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 7650 13920 7656 13932
rect 6549 13883 6607 13889
rect 7576 13892 7656 13920
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2498 13812 2504 13864
rect 2556 13852 2562 13864
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 2556 13824 4537 13852
rect 2556 13812 2562 13824
rect 4525 13821 4537 13824
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4890 13852 4896 13864
rect 4755 13824 4896 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4890 13812 4896 13824
rect 4948 13852 4954 13864
rect 5442 13852 5448 13864
rect 4948 13824 5448 13852
rect 4948 13812 4954 13824
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 5828 13784 5856 13815
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7576 13861 7604 13892
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 11624 13920 11652 14019
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11756 14028 11989 14056
rect 11756 14016 11762 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12345 14059 12403 14065
rect 12345 14056 12357 14059
rect 12124 14028 12357 14056
rect 12124 14016 12130 14028
rect 12345 14025 12357 14028
rect 12391 14025 12403 14059
rect 12345 14019 12403 14025
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 13596 14028 14749 14056
rect 13596 14016 13602 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 17218 14056 17224 14068
rect 15611 14028 17224 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 17368 14028 18889 14056
rect 17368 14016 17374 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 19426 14016 19432 14068
rect 19484 14016 19490 14068
rect 19610 14016 19616 14068
rect 19668 14056 19674 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 19668 14028 20085 14056
rect 19668 14016 19674 14028
rect 20073 14025 20085 14028
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 21232 14028 23397 14056
rect 21232 14016 21238 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 24949 14059 25007 14065
rect 24949 14025 24961 14059
rect 24995 14056 25007 14059
rect 25774 14056 25780 14068
rect 24995 14028 25780 14056
rect 24995 14025 25007 14028
rect 24949 14019 25007 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 11848 13960 13645 13988
rect 11848 13948 11854 13960
rect 13633 13957 13645 13960
rect 13679 13957 13691 13991
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 13633 13951 13691 13957
rect 13740 13960 15945 13988
rect 12066 13920 12072 13932
rect 11624 13892 12072 13920
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 12400 13892 12572 13920
rect 12400 13880 12406 13892
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 7340 13824 7573 13852
rect 7340 13812 7346 13824
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 5902 13784 5908 13796
rect 5828 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 8680 13784 8708 13815
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10100 13824 11069 13852
rect 10100 13812 10106 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 11790 13852 11796 13864
rect 11572 13824 11796 13852
rect 11572 13812 11578 13824
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12544 13861 12572 13892
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 13740 13920 13768 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 16666 13948 16672 14000
rect 16724 13988 16730 14000
rect 17862 13988 17868 14000
rect 16724 13960 17868 13988
rect 16724 13948 16730 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 20990 13948 20996 14000
rect 21048 13988 21054 14000
rect 21048 13960 21772 13988
rect 21048 13948 21054 13960
rect 15194 13920 15200 13932
rect 13648 13892 13768 13920
rect 14752 13892 15200 13920
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12216 13824 12449 13852
rect 12216 13812 12222 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 13648 13852 13676 13892
rect 12860 13824 13676 13852
rect 13817 13855 13875 13861
rect 12860 13812 12866 13824
rect 13817 13821 13829 13855
rect 13863 13821 13875 13855
rect 14752 13852 14780 13892
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16942 13920 16948 13932
rect 16071 13892 16948 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 13817 13815 13875 13821
rect 14384 13824 14780 13852
rect 14829 13855 14887 13861
rect 7708 13756 8708 13784
rect 7708 13744 7714 13756
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 13630 13784 13636 13796
rect 10652 13756 13636 13784
rect 10652 13744 10658 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 5258 13676 5264 13728
rect 5316 13676 5322 13728
rect 5442 13676 5448 13728
rect 5500 13716 5506 13728
rect 5810 13716 5816 13728
rect 5500 13688 5816 13716
rect 5500 13676 5506 13688
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 8938 13716 8944 13728
rect 7524 13688 8944 13716
rect 7524 13676 7530 13688
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 9398 13716 9404 13728
rect 9088 13688 9404 13716
rect 9088 13676 9094 13688
rect 9398 13676 9404 13688
rect 9456 13676 9462 13728
rect 9572 13719 9630 13725
rect 9572 13685 9584 13719
rect 9618 13716 9630 13719
rect 12342 13716 12348 13728
rect 9618 13688 12348 13716
rect 9618 13685 9630 13688
rect 9572 13679 9630 13685
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 13832 13716 13860 13815
rect 14384 13793 14412 13824
rect 14829 13821 14841 13855
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15102 13852 15108 13864
rect 15059 13824 15108 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 14369 13787 14427 13793
rect 14369 13753 14381 13787
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 14844 13784 14872 13815
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 14516 13756 14872 13784
rect 16224 13784 16252 13815
rect 17402 13812 17408 13864
rect 17460 13812 17466 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 19628 13852 19656 13883
rect 20438 13880 20444 13932
rect 20496 13880 20502 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 21634 13920 21640 13932
rect 20579 13892 21640 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 21744 13920 21772 13960
rect 21818 13948 21824 14000
rect 21876 13988 21882 14000
rect 21913 13991 21971 13997
rect 21913 13988 21925 13991
rect 21876 13960 21925 13988
rect 21876 13948 21882 13960
rect 21913 13957 21925 13960
rect 21959 13988 21971 13991
rect 21959 13960 22692 13988
rect 21959 13957 21971 13960
rect 21913 13951 21971 13957
rect 22002 13920 22008 13932
rect 21744 13892 22008 13920
rect 22002 13880 22008 13892
rect 22060 13920 22066 13932
rect 22664 13929 22692 13960
rect 24578 13948 24584 14000
rect 24636 13988 24642 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 24636 13960 25053 13988
rect 24636 13948 24642 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 25314 13948 25320 14000
rect 25372 13988 25378 14000
rect 25593 13991 25651 13997
rect 25593 13988 25605 13991
rect 25372 13960 25605 13988
rect 25372 13948 25378 13960
rect 25593 13957 25605 13960
rect 25639 13957 25651 13991
rect 25593 13951 25651 13957
rect 25682 13948 25688 14000
rect 25740 13988 25746 14000
rect 25869 13991 25927 13997
rect 25869 13988 25881 13991
rect 25740 13960 25881 13988
rect 25740 13948 25746 13960
rect 25869 13957 25881 13960
rect 25915 13957 25927 13991
rect 25869 13951 25927 13957
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22060 13892 22569 13920
rect 22060 13880 22066 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 23753 13923 23811 13929
rect 22695 13892 23244 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 17828 13824 19656 13852
rect 20625 13855 20683 13861
rect 17828 13812 17834 13824
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 20824 13824 22232 13852
rect 20640 13784 20668 13815
rect 20714 13784 20720 13796
rect 16224 13756 17264 13784
rect 20640 13756 20720 13784
rect 14516 13744 14522 13756
rect 16298 13716 16304 13728
rect 13832 13688 16304 13716
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 16666 13676 16672 13728
rect 16724 13676 16730 13728
rect 17236 13716 17264 13756
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 18966 13716 18972 13728
rect 17236 13688 18972 13716
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20824 13716 20852 13824
rect 22204 13793 22232 13824
rect 22189 13787 22247 13793
rect 22189 13753 22201 13787
rect 22235 13753 22247 13787
rect 22572 13784 22600 13883
rect 22830 13812 22836 13864
rect 22888 13812 22894 13864
rect 23216 13852 23244 13892
rect 23753 13889 23765 13923
rect 23799 13920 23811 13923
rect 25961 13923 26019 13929
rect 25961 13920 25973 13923
rect 23799 13892 25973 13920
rect 23799 13889 23811 13892
rect 23753 13883 23811 13889
rect 23842 13852 23848 13864
rect 23216 13824 23848 13852
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 23952 13784 23980 13892
rect 25961 13889 25973 13892
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 24026 13812 24032 13864
rect 24084 13812 24090 13864
rect 25133 13855 25191 13861
rect 25133 13821 25145 13855
rect 25179 13821 25191 13855
rect 25133 13815 25191 13821
rect 22572 13756 23980 13784
rect 22189 13747 22247 13753
rect 24118 13744 24124 13796
rect 24176 13784 24182 13796
rect 25148 13784 25176 13815
rect 24176 13756 25176 13784
rect 24176 13744 24182 13756
rect 20220 13688 20852 13716
rect 20220 13676 20226 13688
rect 21910 13676 21916 13728
rect 21968 13716 21974 13728
rect 22554 13716 22560 13728
rect 21968 13688 22560 13716
rect 21968 13676 21974 13688
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 24578 13676 24584 13728
rect 24636 13676 24642 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 5224 13484 5672 13512
rect 5224 13472 5230 13484
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13376 4215 13379
rect 5166 13376 5172 13388
rect 4203 13348 5172 13376
rect 4203 13345 4215 13348
rect 4157 13339 4215 13345
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5644 13376 5672 13484
rect 6270 13472 6276 13524
rect 6328 13472 6334 13524
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 10134 13512 10140 13524
rect 7800 13484 10140 13512
rect 7800 13472 7806 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 10744 13484 11621 13512
rect 10744 13472 10750 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 10594 13444 10600 13456
rect 9140 13416 10600 13444
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 5644 13348 6745 13376
rect 6733 13345 6745 13348
rect 6779 13376 6791 13379
rect 7374 13376 7380 13388
rect 6779 13348 7380 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 9030 13376 9036 13388
rect 7800 13348 9036 13376
rect 7800 13336 7806 13348
rect 9030 13336 9036 13348
rect 9088 13336 9094 13388
rect 9140 13385 9168 13416
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11425 13447 11483 13453
rect 11425 13444 11437 13447
rect 11112 13416 11437 13444
rect 11112 13404 11118 13416
rect 11425 13413 11437 13416
rect 11471 13413 11483 13447
rect 11425 13407 11483 13413
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 6270 13308 6276 13320
rect 5566 13280 6276 13308
rect 1765 13271 1823 13277
rect 1780 13240 1808 13271
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 10980 13308 11008 13339
rect 8496 13280 11008 13308
rect 3326 13240 3332 13252
rect 1780 13212 3332 13240
rect 3326 13200 3332 13212
rect 3384 13200 3390 13252
rect 4430 13200 4436 13252
rect 4488 13200 4494 13252
rect 6914 13240 6920 13252
rect 5736 13212 6920 13240
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 5736 13172 5764 13212
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7282 13240 7288 13252
rect 7055 13212 7288 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7392 13212 7498 13240
rect 1912 13144 5764 13172
rect 1912 13132 1918 13144
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6270 13132 6276 13184
rect 6328 13172 6334 13184
rect 7392 13172 7420 13212
rect 6328 13144 7420 13172
rect 6328 13132 6334 13144
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8496 13181 8524 13280
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 9582 13240 9588 13252
rect 8812 13212 9588 13240
rect 8812 13200 8818 13212
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 10873 13243 10931 13249
rect 10873 13240 10885 13243
rect 9732 13212 10885 13240
rect 9732 13200 9738 13212
rect 10873 13209 10885 13212
rect 10919 13209 10931 13243
rect 10873 13203 10931 13209
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 7708 13144 8493 13172
rect 7708 13132 7714 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 9490 13132 9496 13184
rect 9548 13172 9554 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9548 13144 10425 13172
rect 9548 13132 9554 13144
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10413 13135 10471 13141
rect 10778 13132 10784 13184
rect 10836 13132 10842 13184
rect 11624 13172 11652 13475
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 12308 13484 13737 13512
rect 12308 13472 12314 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15068 13484 16037 13512
rect 15068 13472 15074 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 17460 13484 18889 13512
rect 17460 13472 17466 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 21910 13512 21916 13524
rect 18877 13475 18935 13481
rect 18984 13484 21916 13512
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 18984 13444 19012 13484
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22646 13512 22652 13524
rect 22143 13484 22652 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23937 13515 23995 13521
rect 23937 13512 23949 13515
rect 23164 13484 23949 13512
rect 23164 13472 23170 13484
rect 23937 13481 23949 13484
rect 23983 13512 23995 13515
rect 24486 13512 24492 13524
rect 23983 13484 24492 13512
rect 23983 13481 23995 13484
rect 23937 13475 23995 13481
rect 24486 13472 24492 13484
rect 24544 13472 24550 13524
rect 18840 13416 19012 13444
rect 18840 13404 18846 13416
rect 21634 13404 21640 13456
rect 21692 13444 21698 13456
rect 22833 13447 22891 13453
rect 22833 13444 22845 13447
rect 21692 13416 22845 13444
rect 21692 13404 21698 13416
rect 22833 13413 22845 13416
rect 22879 13413 22891 13447
rect 23750 13444 23756 13456
rect 22833 13407 22891 13413
rect 23308 13416 23756 13444
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 13262 13376 13268 13388
rect 12032 13348 13268 13376
rect 12032 13336 12038 13348
rect 13262 13336 13268 13348
rect 13320 13376 13326 13388
rect 14553 13379 14611 13385
rect 13320 13348 14320 13376
rect 13320 13336 13326 13348
rect 14292 13320 14320 13348
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15194 13376 15200 13388
rect 14599 13348 15200 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15194 13336 15200 13348
rect 15252 13376 15258 13388
rect 16390 13376 16396 13388
rect 15252 13348 16396 13376
rect 15252 13336 15258 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 17126 13336 17132 13388
rect 17184 13336 17190 13388
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 20349 13379 20407 13385
rect 17920 13348 18552 13376
rect 17920 13336 17926 13348
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 12250 13200 12256 13252
rect 12308 13200 12314 13252
rect 12710 13240 12716 13252
rect 12636 13212 12716 13240
rect 12636 13172 12664 13212
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14240 13212 15042 13240
rect 14240 13200 14246 13212
rect 16298 13200 16304 13252
rect 16356 13240 16362 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 16356 13212 17417 13240
rect 16356 13200 16362 13212
rect 17405 13209 17417 13212
rect 17451 13209 17463 13243
rect 17405 13203 17463 13209
rect 11624 13144 12664 13172
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 16485 13175 16543 13181
rect 16485 13172 16497 13175
rect 14700 13144 16497 13172
rect 14700 13132 14706 13144
rect 16485 13141 16497 13144
rect 16531 13141 16543 13175
rect 17420 13172 17448 13203
rect 17862 13200 17868 13252
rect 17920 13200 17926 13252
rect 18322 13172 18328 13184
rect 17420 13144 18328 13172
rect 16485 13135 16543 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18524 13172 18552 13348
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 22186 13376 22192 13388
rect 20395 13348 22192 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 23308 13385 23336 13416
rect 23750 13404 23756 13416
rect 23808 13404 23814 13456
rect 23842 13404 23848 13456
rect 23900 13444 23906 13456
rect 24121 13447 24179 13453
rect 24121 13444 24133 13447
rect 23900 13416 24133 13444
rect 23900 13404 23906 13416
rect 24121 13413 24133 13416
rect 24167 13413 24179 13447
rect 24121 13407 24179 13413
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 23474 13336 23480 13388
rect 23532 13336 23538 13388
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 32490 13376 32496 13388
rect 23624 13348 32496 13376
rect 23624 13336 23630 13348
rect 32490 13336 32496 13348
rect 32548 13336 32554 13388
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 22002 13268 22008 13320
rect 22060 13308 22066 13320
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22060 13280 22477 13308
rect 22060 13268 22066 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23072 13280 25452 13308
rect 23072 13268 23078 13280
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 19024 13212 20637 13240
rect 19024 13200 19030 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 23201 13243 23259 13249
rect 23201 13209 23213 13243
rect 23247 13240 23259 13243
rect 23247 13212 23336 13240
rect 23247 13209 23259 13212
rect 23201 13203 23259 13209
rect 19337 13175 19395 13181
rect 19337 13172 19349 13175
rect 18524 13144 19349 13172
rect 19337 13141 19349 13144
rect 19383 13172 19395 13175
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 19383 13144 19441 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 22922 13172 22928 13184
rect 20404 13144 22928 13172
rect 20404 13132 20410 13144
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 23308 13172 23336 13212
rect 24486 13200 24492 13252
rect 24544 13240 24550 13252
rect 25424 13249 25452 13280
rect 24581 13243 24639 13249
rect 24581 13240 24593 13243
rect 24544 13212 24593 13240
rect 24544 13200 24550 13212
rect 24581 13209 24593 13212
rect 24627 13209 24639 13243
rect 24581 13203 24639 13209
rect 25409 13243 25467 13249
rect 25409 13209 25421 13243
rect 25455 13240 25467 13243
rect 29730 13240 29736 13252
rect 25455 13212 29736 13240
rect 25455 13209 25467 13212
rect 25409 13203 25467 13209
rect 29730 13200 29736 13212
rect 29788 13200 29794 13252
rect 25222 13172 25228 13184
rect 23308 13144 25228 13172
rect 25222 13132 25228 13144
rect 25280 13132 25286 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 4982 12928 4988 12980
rect 5040 12928 5046 12980
rect 5718 12928 5724 12980
rect 5776 12928 5782 12980
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 7098 12968 7104 12980
rect 6604 12940 7104 12968
rect 6604 12928 6610 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 9858 12968 9864 12980
rect 7331 12940 9864 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 10505 12971 10563 12977
rect 10505 12968 10517 12971
rect 10192 12940 10517 12968
rect 10192 12928 10198 12940
rect 10505 12937 10517 12940
rect 10551 12937 10563 12971
rect 10505 12931 10563 12937
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10744 12940 10977 12968
rect 10744 12928 10750 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 11204 12940 12541 12968
rect 11204 12928 11210 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 15378 12968 15384 12980
rect 12529 12931 12587 12937
rect 13096 12940 15384 12968
rect 3694 12860 3700 12912
rect 3752 12860 3758 12912
rect 4249 12903 4307 12909
rect 4249 12869 4261 12903
rect 4295 12900 4307 12903
rect 4338 12900 4344 12912
rect 4295 12872 4344 12900
rect 4295 12869 4307 12872
rect 4249 12863 4307 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 5629 12903 5687 12909
rect 5629 12869 5641 12903
rect 5675 12900 5687 12903
rect 5810 12900 5816 12912
rect 5675 12872 5816 12900
rect 5675 12869 5687 12872
rect 5629 12863 5687 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 8570 12900 8576 12912
rect 7064 12872 8576 12900
rect 7064 12860 7070 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 8754 12860 8760 12912
rect 8812 12860 8818 12912
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 10704 12900 10732 12928
rect 9640 12872 10732 12900
rect 11885 12903 11943 12909
rect 9640 12860 9646 12872
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 12434 12900 12440 12912
rect 11931 12872 12440 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1360 12804 1593 12832
rect 1360 12792 1366 12804
rect 1581 12801 1593 12804
rect 1627 12832 1639 12835
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 1627 12804 2697 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 3786 12832 3792 12844
rect 3559 12804 3792 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 4488 12804 5948 12832
rect 4488 12792 4494 12804
rect 1854 12724 1860 12776
rect 1912 12724 1918 12776
rect 3418 12724 3424 12776
rect 3476 12764 3482 12776
rect 3694 12764 3700 12776
rect 3476 12736 3700 12764
rect 3476 12724 3482 12736
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 5920 12773 5948 12804
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 6972 12804 7205 12832
rect 6972 12792 6978 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 10318 12832 10324 12844
rect 10091 12804 10324 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12406 12804 12909 12832
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 5951 12736 7389 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 9030 12764 9036 12776
rect 8343 12736 9036 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 4433 12699 4491 12705
rect 4433 12665 4445 12699
rect 4479 12696 4491 12699
rect 7742 12696 7748 12708
rect 4479 12668 7748 12696
rect 4479 12665 4491 12668
rect 4433 12659 4491 12665
rect 7742 12656 7748 12668
rect 7800 12656 7806 12708
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5626 12628 5632 12640
rect 5307 12600 5632 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 6822 12588 6828 12640
rect 6880 12588 6886 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 8036 12628 8064 12727
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 12406 12764 12434 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 10192 12736 12434 12764
rect 10192 12724 10198 12736
rect 12986 12724 12992 12776
rect 13044 12724 13050 12776
rect 13096 12773 13124 12940
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17000 12940 17785 12968
rect 17000 12928 17006 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 20162 12968 20168 12980
rect 18187 12940 20168 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21174 12968 21180 12980
rect 21131 12940 21180 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21726 12928 21732 12980
rect 21784 12968 21790 12980
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 21784 12940 22201 12968
rect 21784 12928 21790 12940
rect 22189 12937 22201 12940
rect 22235 12937 22247 12971
rect 22189 12931 22247 12937
rect 22922 12928 22928 12980
rect 22980 12968 22986 12980
rect 23474 12968 23480 12980
rect 22980 12940 23480 12968
rect 22980 12928 22986 12940
rect 23474 12928 23480 12940
rect 23532 12968 23538 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23532 12940 24777 12968
rect 23532 12928 23538 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 14093 12903 14151 12909
rect 14093 12900 14105 12903
rect 14016 12872 14105 12900
rect 13262 12792 13268 12844
rect 13320 12832 13326 12844
rect 14016 12832 14044 12872
rect 14093 12869 14105 12872
rect 14139 12869 14151 12903
rect 14093 12863 14151 12869
rect 14274 12860 14280 12912
rect 14332 12900 14338 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 14332 12872 15669 12900
rect 14332 12860 14338 12872
rect 15657 12869 15669 12872
rect 15703 12869 15715 12903
rect 15657 12863 15715 12869
rect 16393 12903 16451 12909
rect 16393 12869 16405 12903
rect 16439 12900 16451 12903
rect 18414 12900 18420 12912
rect 16439 12872 18420 12900
rect 16439 12869 16451 12872
rect 16393 12863 16451 12869
rect 13320 12804 14044 12832
rect 13320 12792 13326 12804
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 16408 12832 16436 12863
rect 18414 12860 18420 12872
rect 18472 12900 18478 12912
rect 18874 12900 18880 12912
rect 18472 12872 18880 12900
rect 18472 12860 18478 12872
rect 18874 12860 18880 12872
rect 18932 12900 18938 12912
rect 18969 12903 19027 12909
rect 18969 12900 18981 12903
rect 18932 12872 18981 12900
rect 18932 12860 18938 12872
rect 18969 12869 18981 12872
rect 19015 12869 19027 12903
rect 18969 12863 19027 12869
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 23566 12900 23572 12912
rect 19208 12872 23572 12900
rect 19208 12860 19214 12872
rect 23566 12860 23572 12872
rect 23624 12860 23630 12912
rect 23934 12860 23940 12912
rect 23992 12860 23998 12912
rect 14976 12804 16436 12832
rect 18233 12835 18291 12841
rect 14976 12792 14982 12804
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 18690 12832 18696 12844
rect 18279 12804 18696 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12832 21235 12835
rect 21542 12832 21548 12844
rect 21223 12804 21548 12832
rect 21223 12801 21235 12804
rect 21177 12795 21235 12801
rect 21542 12792 21548 12804
rect 21600 12792 21606 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23014 12832 23020 12844
rect 22244 12804 23020 12832
rect 22244 12792 22250 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12764 14243 12767
rect 14274 12764 14280 12776
rect 14231 12736 14280 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 15102 12764 15108 12776
rect 14415 12736 15108 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15252 12736 16865 12764
rect 15252 12724 15258 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 18414 12724 18420 12776
rect 18472 12724 18478 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20070 12764 20076 12776
rect 19843 12736 20076 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12696 11299 12699
rect 14918 12696 14924 12708
rect 11287 12668 14924 12696
rect 11287 12665 11299 12668
rect 11241 12659 11299 12665
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 18506 12656 18512 12708
rect 18564 12696 18570 12708
rect 19812 12696 19840 12727
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 24302 12764 24308 12776
rect 23339 12736 24308 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 24302 12724 24308 12736
rect 24360 12724 24366 12776
rect 22462 12696 22468 12708
rect 18564 12668 19840 12696
rect 20640 12668 22468 12696
rect 18564 12656 18570 12668
rect 9306 12628 9312 12640
rect 7432 12600 9312 12628
rect 7432 12588 7438 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 11606 12588 11612 12640
rect 11664 12588 11670 12640
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 13262 12628 13268 12640
rect 12216 12600 13268 12628
rect 12216 12588 12222 12600
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 13725 12631 13783 12637
rect 13725 12597 13737 12631
rect 13771 12628 13783 12631
rect 14550 12628 14556 12640
rect 13771 12600 14556 12628
rect 13771 12597 13783 12600
rect 13725 12591 13783 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15344 12600 16129 12628
rect 15344 12588 15350 12600
rect 16117 12597 16129 12600
rect 16163 12628 16175 12631
rect 16666 12628 16672 12640
rect 16163 12600 16672 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 16666 12588 16672 12600
rect 16724 12628 16730 12640
rect 17034 12628 17040 12640
rect 16724 12600 17040 12628
rect 16724 12588 16730 12600
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 20640 12628 20668 12668
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 18748 12600 20668 12628
rect 20717 12631 20775 12637
rect 18748 12588 18754 12600
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 20898 12628 20904 12640
rect 20763 12600 20904 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 23934 12588 23940 12640
rect 23992 12628 23998 12640
rect 24394 12628 24400 12640
rect 23992 12600 24400 12628
rect 23992 12588 23998 12600
rect 24394 12588 24400 12600
rect 24452 12628 24458 12640
rect 25041 12631 25099 12637
rect 25041 12628 25053 12631
rect 24452 12600 25053 12628
rect 24452 12588 24458 12600
rect 25041 12597 25053 12600
rect 25087 12597 25099 12631
rect 25041 12591 25099 12597
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 2924 12396 3065 12424
rect 2924 12384 2930 12396
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 3053 12387 3111 12393
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4338 12424 4344 12436
rect 4019 12396 4344 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 4706 12424 4712 12436
rect 4663 12396 4712 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 9674 12424 9680 12436
rect 7883 12396 9680 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11793 12427 11851 12433
rect 10980 12396 11744 12424
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 4522 12288 4528 12300
rect 1903 12260 4528 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 4724 12297 4752 12384
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 7340 12328 7880 12356
rect 7340 12316 7346 12328
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5224 12260 5365 12288
rect 5224 12248 5230 12260
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 7742 12288 7748 12300
rect 7423 12260 7748 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 7852 12288 7880 12328
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 10980 12356 11008 12396
rect 11606 12356 11612 12368
rect 8260 12328 11008 12356
rect 11072 12328 11612 12356
rect 8260 12316 8266 12328
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7852 12260 8401 12288
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9364 12260 9873 12288
rect 9364 12248 9370 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1360 12192 1593 12220
rect 1360 12180 1366 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 3007 12192 3433 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3421 12189 3433 12192
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 4154 12220 4160 12232
rect 3927 12192 4160 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 2498 12152 2504 12164
rect 2004 12124 2504 12152
rect 2004 12112 2010 12124
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 3436 12152 3464 12183
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4798 12220 4804 12232
rect 4396 12192 4804 12220
rect 4396 12180 4402 12192
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 8202 12220 8208 12232
rect 7524 12192 8208 12220
rect 7524 12180 7530 12192
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 10410 12220 10416 12232
rect 8343 12192 10416 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11072 12229 11100 12328
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 11238 12248 11244 12300
rect 11296 12248 11302 12300
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12189 11115 12223
rect 11716 12220 11744 12396
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 12526 12424 12532 12436
rect 11839 12396 12532 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 14182 12384 14188 12436
rect 14240 12384 14246 12436
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14332 12396 14381 12424
rect 14332 12384 14338 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14476 12396 17632 12424
rect 14090 12356 14096 12368
rect 11808 12328 14096 12356
rect 11808 12300 11836 12328
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 14476 12356 14504 12396
rect 14200 12328 14504 12356
rect 17604 12356 17632 12396
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18782 12424 18788 12436
rect 18104 12396 18788 12424
rect 18104 12384 18110 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21821 12427 21879 12433
rect 21821 12424 21833 12427
rect 20772 12396 21833 12424
rect 20772 12384 20778 12396
rect 21821 12393 21833 12396
rect 21867 12424 21879 12427
rect 21867 12396 22094 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 19886 12356 19892 12368
rect 17604 12328 19892 12356
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 12345 12291 12403 12297
rect 12345 12288 12357 12291
rect 12308 12260 12357 12288
rect 12308 12248 12314 12260
rect 12345 12257 12357 12260
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 14200 12288 14228 12328
rect 19886 12316 19892 12328
rect 19944 12316 19950 12368
rect 15194 12288 15200 12300
rect 13679 12260 14228 12288
rect 14292 12260 15200 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 11716 12192 12173 12220
rect 11057 12183 11115 12189
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 14292 12220 14320 12260
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 16206 12288 16212 12300
rect 15436 12260 16212 12288
rect 15436 12248 15442 12260
rect 16206 12248 16212 12260
rect 16264 12288 16270 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16264 12260 16589 12288
rect 16264 12248 16270 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 18322 12288 18328 12300
rect 17092 12260 18328 12288
rect 17092 12248 17098 12260
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 20346 12248 20352 12300
rect 20404 12248 20410 12300
rect 22066 12288 22094 12396
rect 24394 12384 24400 12436
rect 24452 12384 24458 12436
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 22066 12260 22569 12288
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 13403 12192 14320 12220
rect 14737 12223 14795 12229
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14918 12220 14924 12232
rect 14783 12192 14924 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14918 12180 14924 12192
rect 14976 12220 14982 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 14976 12192 15945 12220
rect 14976 12180 14982 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 16301 12183 16359 12189
rect 17972 12192 19533 12220
rect 5534 12152 5540 12164
rect 3436 12124 5540 12152
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 5629 12155 5687 12161
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5718 12152 5724 12164
rect 5675 12124 5724 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 6270 12112 6276 12164
rect 6328 12112 6334 12164
rect 9122 12112 9128 12164
rect 9180 12152 9186 12164
rect 9950 12152 9956 12164
rect 9180 12124 9956 12152
rect 9180 12112 9186 12124
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 10060 12124 14412 12152
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 6972 12056 8217 12084
rect 6972 12044 6978 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 10060 12084 10088 12124
rect 8996 12056 10088 12084
rect 8996 12044 9002 12056
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 10744 12056 10977 12084
rect 10744 12044 10750 12056
rect 10965 12053 10977 12056
rect 11011 12053 11023 12087
rect 10965 12047 11023 12053
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 12066 12084 12072 12096
rect 11296 12056 12072 12084
rect 11296 12044 11302 12056
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12250 12044 12256 12096
rect 12308 12044 12314 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13262 12084 13268 12096
rect 13035 12056 13268 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 13446 12044 13452 12096
rect 13504 12044 13510 12096
rect 14384 12084 14412 12124
rect 14458 12112 14464 12164
rect 14516 12152 14522 12164
rect 15473 12155 15531 12161
rect 15473 12152 15485 12155
rect 14516 12124 15485 12152
rect 14516 12112 14522 12124
rect 15473 12121 15485 12124
rect 15519 12152 15531 12155
rect 16316 12152 16344 12183
rect 15519 12124 16344 12152
rect 15519 12121 15531 12124
rect 15473 12115 15531 12121
rect 17034 12112 17040 12164
rect 17092 12112 17098 12164
rect 17402 12084 17408 12096
rect 14384 12056 17408 12084
rect 17402 12044 17408 12056
rect 17460 12084 17466 12096
rect 17972 12084 18000 12192
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 18322 12112 18328 12164
rect 18380 12152 18386 12164
rect 18380 12124 18644 12152
rect 18380 12112 18386 12124
rect 17460 12056 18000 12084
rect 17460 12044 17466 12056
rect 18506 12044 18512 12096
rect 18564 12044 18570 12096
rect 18616 12084 18644 12124
rect 18874 12112 18880 12164
rect 18932 12152 18938 12164
rect 18932 12124 19288 12152
rect 18932 12112 18938 12124
rect 19260 12096 19288 12124
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18616 12056 18981 12084
rect 18969 12053 18981 12056
rect 19015 12053 19027 12087
rect 18969 12047 19027 12053
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 19300 12056 19349 12084
rect 19300 12044 19306 12056
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19536 12084 19564 12183
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22244 12192 22293 12220
rect 22244 12180 22250 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 23934 12220 23940 12232
rect 23690 12192 23940 12220
rect 22281 12183 22339 12189
rect 23934 12180 23940 12192
rect 23992 12180 23998 12232
rect 21726 12152 21732 12164
rect 21574 12124 21732 12152
rect 21726 12112 21732 12124
rect 21784 12112 21790 12164
rect 25038 12152 25044 12164
rect 23952 12124 25044 12152
rect 23952 12084 23980 12124
rect 25038 12112 25044 12124
rect 25096 12112 25102 12164
rect 19536 12056 23980 12084
rect 19337 12047 19395 12053
rect 24026 12044 24032 12096
rect 24084 12044 24090 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1302 11840 1308 11892
rect 1360 11880 1366 11892
rect 1397 11883 1455 11889
rect 1397 11880 1409 11883
rect 1360 11852 1409 11880
rect 1360 11840 1366 11852
rect 1397 11849 1409 11852
rect 1443 11849 1455 11883
rect 1397 11843 1455 11849
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4479 11852 5273 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 11701 11883 11759 11889
rect 6779 11852 10088 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 3329 11815 3387 11821
rect 3329 11781 3341 11815
rect 3375 11812 3387 11815
rect 3421 11815 3479 11821
rect 3421 11812 3433 11815
rect 3375 11784 3433 11812
rect 3375 11781 3387 11784
rect 3329 11775 3387 11781
rect 3421 11781 3433 11784
rect 3467 11812 3479 11815
rect 5721 11815 5779 11821
rect 3467 11784 5396 11812
rect 3467 11781 3479 11784
rect 3421 11775 3479 11781
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 2372 11716 2421 11744
rect 2372 11704 2378 11716
rect 2409 11713 2421 11716
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 5258 11744 5264 11756
rect 4571 11716 5264 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5368 11744 5396 11784
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6822 11812 6828 11824
rect 5767 11784 6828 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7650 11772 7656 11824
rect 7708 11772 7714 11824
rect 8202 11772 8208 11824
rect 8260 11772 8266 11824
rect 6546 11744 6552 11756
rect 5368 11716 6552 11744
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 9950 11744 9956 11756
rect 9631 11716 9956 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10060 11744 10088 11852
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 12250 11880 12256 11892
rect 11747 11852 12256 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 12250 11840 12256 11852
rect 12308 11880 12314 11892
rect 12802 11880 12808 11892
rect 12308 11852 12808 11880
rect 12308 11840 12314 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 15194 11840 15200 11892
rect 15252 11840 15258 11892
rect 15562 11840 15568 11892
rect 15620 11840 15626 11892
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 16071 11852 17356 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 12437 11815 12495 11821
rect 12437 11812 12449 11815
rect 10652 11784 12449 11812
rect 10652 11772 10658 11784
rect 12437 11781 12449 11784
rect 12483 11781 12495 11815
rect 13354 11812 13360 11824
rect 12437 11775 12495 11781
rect 13188 11784 13360 11812
rect 13188 11753 13216 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 14182 11772 14188 11824
rect 14240 11772 14246 11824
rect 17328 11812 17356 11852
rect 17402 11840 17408 11892
rect 17460 11840 17466 11892
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 18141 11883 18199 11889
rect 18141 11880 18153 11883
rect 17828 11852 18153 11880
rect 17828 11840 17834 11852
rect 18141 11849 18153 11852
rect 18187 11849 18199 11883
rect 18141 11843 18199 11849
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 19337 11883 19395 11889
rect 19337 11880 19349 11883
rect 18656 11852 19349 11880
rect 18656 11840 18662 11852
rect 19337 11849 19349 11852
rect 19383 11849 19395 11883
rect 20898 11880 20904 11892
rect 19337 11843 19395 11849
rect 19444 11852 20904 11880
rect 17328 11784 17540 11812
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 10060 11716 12357 11744
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 14792 11716 15945 11744
rect 14792 11704 14798 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 16172 11716 17325 11744
rect 16172 11704 16178 11716
rect 17313 11713 17325 11716
rect 17359 11713 17371 11747
rect 17512 11744 17540 11784
rect 17586 11772 17592 11824
rect 17644 11812 17650 11824
rect 18509 11815 18567 11821
rect 18509 11812 18521 11815
rect 17644 11784 18521 11812
rect 17644 11772 17650 11784
rect 18509 11781 18521 11784
rect 18555 11812 18567 11815
rect 19153 11815 19211 11821
rect 19153 11812 19165 11815
rect 18555 11784 19165 11812
rect 18555 11781 18567 11784
rect 18509 11775 18567 11781
rect 19153 11781 19165 11784
rect 19199 11781 19211 11815
rect 19153 11775 19211 11781
rect 19444 11744 19472 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21726 11840 21732 11892
rect 21784 11880 21790 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 21784 11852 21925 11880
rect 21784 11840 21790 11852
rect 21913 11849 21925 11852
rect 21959 11849 21971 11883
rect 24026 11880 24032 11892
rect 21913 11843 21971 11849
rect 22112 11852 24032 11880
rect 21744 11812 21772 11840
rect 21206 11784 21772 11812
rect 17512 11716 19472 11744
rect 17313 11707 17371 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2130 11676 2136 11688
rect 2004 11648 2136 11676
rect 2004 11636 2010 11648
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 4062 11676 4068 11688
rect 2832 11648 4068 11676
rect 2832 11636 2838 11648
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 5626 11676 5632 11688
rect 4755 11648 5632 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5902 11636 5908 11688
rect 5960 11636 5966 11688
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 8110 11676 8116 11688
rect 7248 11648 8116 11676
rect 7248 11636 7254 11648
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 8680 11648 10333 11676
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5920 11608 5948 11636
rect 5592 11580 5948 11608
rect 5592 11568 5598 11580
rect 7006 11568 7012 11620
rect 7064 11608 7070 11620
rect 7374 11608 7380 11620
rect 7064 11580 7380 11608
rect 7064 11568 7070 11580
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 7650 11540 7656 11552
rect 4111 11512 7656 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8680 11540 8708 11648
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 11790 11676 11796 11688
rect 11011 11648 11796 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 9030 11568 9036 11620
rect 9088 11608 9094 11620
rect 9125 11611 9183 11617
rect 9125 11608 9137 11611
rect 9088 11580 9137 11608
rect 9088 11568 9094 11580
rect 9125 11577 9137 11580
rect 9171 11577 9183 11611
rect 10336 11608 10364 11639
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 12250 11636 12256 11688
rect 12308 11676 12314 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12308 11648 12541 11676
rect 12308 11636 12314 11648
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 15010 11676 15016 11688
rect 13495 11648 15016 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 17034 11676 17040 11688
rect 16255 11648 17040 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 11514 11608 11520 11620
rect 10336 11580 11520 11608
rect 9125 11571 9183 11577
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 17328 11608 17356 11707
rect 17586 11636 17592 11688
rect 17644 11636 17650 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18616 11648 18705 11676
rect 18506 11608 18512 11620
rect 15028 11580 17264 11608
rect 17328 11580 18512 11608
rect 15028 11552 15056 11580
rect 7892 11512 8708 11540
rect 7892 11500 7898 11512
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 10502 11540 10508 11552
rect 8812 11512 10508 11540
rect 8812 11500 8818 11512
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 12124 11512 14933 11540
rect 12124 11500 12130 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 15010 11500 15016 11552
rect 15068 11500 15074 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 15344 11512 16957 11540
rect 15344 11500 15350 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 17236 11540 17264 11580
rect 18506 11568 18512 11580
rect 18564 11568 18570 11620
rect 18616 11540 18644 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 19702 11636 19708 11688
rect 19760 11636 19766 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11676 20039 11679
rect 22112 11676 22140 11852
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 24394 11840 24400 11892
rect 24452 11840 24458 11892
rect 22649 11815 22707 11821
rect 22649 11781 22661 11815
rect 22695 11812 22707 11815
rect 22738 11812 22744 11824
rect 22695 11784 22744 11812
rect 22695 11781 22707 11784
rect 22649 11775 22707 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 23934 11812 23940 11824
rect 23874 11784 23940 11812
rect 23934 11772 23940 11784
rect 23992 11812 23998 11824
rect 24412 11812 24440 11840
rect 23992 11784 24440 11812
rect 23992 11772 23998 11784
rect 20027 11648 22140 11676
rect 20027 11645 20039 11648
rect 19981 11639 20039 11645
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22244 11648 22385 11676
rect 22244 11636 22250 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 17236 11512 18644 11540
rect 16945 11503 17003 11509
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 24118 11500 24124 11552
rect 24176 11500 24182 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 2240 11308 3280 11336
rect 2240 11209 2268 11308
rect 2774 11268 2780 11280
rect 2332 11240 2780 11268
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2332 11132 2360 11240
rect 2774 11228 2780 11240
rect 2832 11228 2838 11280
rect 2498 11160 2504 11212
rect 2556 11160 2562 11212
rect 3252 11200 3280 11308
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 3602 11336 3608 11348
rect 3476 11308 3608 11336
rect 3476 11296 3482 11308
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 5064 11339 5122 11345
rect 5064 11305 5076 11339
rect 5110 11336 5122 11339
rect 5534 11336 5540 11348
rect 5110 11308 5540 11336
rect 5110 11305 5122 11308
rect 5064 11299 5122 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5776 11308 6561 11336
rect 5776 11296 5782 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 12526 11336 12532 11348
rect 6549 11299 6607 11305
rect 6932 11308 12532 11336
rect 4246 11228 4252 11280
rect 4304 11228 4310 11280
rect 3252 11172 3464 11200
rect 3436 11141 3464 11172
rect 3602 11160 3608 11212
rect 3660 11160 3666 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 6822 11200 6828 11212
rect 4847 11172 6828 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 1811 11104 2360 11132
rect 3421 11135 3479 11141
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 6362 11132 6368 11144
rect 3467 11104 4844 11132
rect 6210 11104 6368 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 1596 11036 4077 11064
rect 1596 11005 1624 11036
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4816 11064 4844 11104
rect 6362 11092 6368 11104
rect 6420 11132 6426 11144
rect 6730 11132 6736 11144
rect 6420 11104 6736 11132
rect 6420 11092 6426 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6932 11064 6960 11308
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 13504 11308 13645 11336
rect 13504 11296 13510 11308
rect 13633 11305 13645 11308
rect 13679 11336 13691 11339
rect 14182 11336 14188 11348
rect 13679 11308 14188 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 16114 11336 16120 11348
rect 14844 11308 16120 11336
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 7800 11240 7849 11268
rect 7800 11228 7806 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 8754 11268 8760 11280
rect 7837 11231 7895 11237
rect 7944 11240 8760 11268
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7944 11132 7972 11240
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9088 11240 9720 11268
rect 9088 11228 9094 11240
rect 8110 11160 8116 11212
rect 8168 11200 8174 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8168 11172 8401 11200
rect 8168 11160 8174 11172
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 9692 11209 9720 11240
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 14844 11268 14872 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 16264 11308 16497 11336
rect 16264 11296 16270 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 18966 11336 18972 11348
rect 18923 11308 18972 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 22830 11336 22836 11348
rect 22695 11308 22836 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23017 11339 23075 11345
rect 23017 11305 23029 11339
rect 23063 11336 23075 11339
rect 23934 11336 23940 11348
rect 23063 11308 23940 11336
rect 23063 11305 23075 11308
rect 23017 11299 23075 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 30098 11296 30104 11348
rect 30156 11336 30162 11348
rect 32033 11339 32091 11345
rect 32033 11336 32045 11339
rect 30156 11308 32045 11336
rect 30156 11296 30162 11308
rect 32033 11305 32045 11308
rect 32079 11305 32091 11339
rect 32033 11299 32091 11305
rect 12860 11240 14872 11268
rect 12860 11228 12866 11240
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9272 11172 9597 11200
rect 9272 11160 9278 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10226 11200 10232 11212
rect 9824 11172 10232 11200
rect 9824 11160 9830 11172
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 7055 11104 7972 11132
rect 8205 11135 8263 11141
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8294 11132 8300 11144
rect 8251 11104 8300 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 4816 11036 5488 11064
rect 4065 11027 4123 11033
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10965 1639 10999
rect 5460 10996 5488 11036
rect 6380 11036 6960 11064
rect 6380 10996 6408 11036
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 7984 11036 8340 11064
rect 7984 11024 7990 11036
rect 5460 10968 6408 10996
rect 1581 10959 1639 10965
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 7469 10999 7527 11005
rect 7469 10996 7481 10999
rect 6788 10968 7481 10996
rect 6788 10956 6794 10968
rect 7469 10965 7481 10968
rect 7515 10996 7527 10999
rect 8202 10996 8208 11008
rect 7515 10968 8208 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8312 11005 8340 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 9456 11036 10701 11064
rect 9456 11024 9462 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10980 11064 11008 11163
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 12400 11172 13277 11200
rect 12400 11160 12406 11172
rect 13265 11169 13277 11172
rect 13311 11169 13323 11203
rect 13265 11163 13323 11169
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 19978 11200 19984 11212
rect 13412 11172 19984 11200
rect 13412 11160 13418 11172
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 29730 11160 29736 11212
rect 29788 11160 29794 11212
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14516 11104 14749 11132
rect 14516 11092 14522 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16908 11104 17141 11132
rect 16908 11092 16914 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 19242 11092 19248 11144
rect 19300 11132 19306 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 19300 11104 19533 11132
rect 19300 11092 19306 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 10980 11036 11805 11064
rect 10689 11027 10747 11033
rect 11793 11033 11805 11036
rect 11839 11064 11851 11067
rect 13446 11064 13452 11076
rect 11839 11036 12204 11064
rect 13018 11036 13452 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10965 8355 10999
rect 8297 10959 8355 10965
rect 9125 10999 9183 11005
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 9214 10996 9220 11008
rect 9171 10968 9220 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 10318 10956 10324 11008
rect 10376 10956 10382 11008
rect 10778 10956 10784 11008
rect 10836 10956 10842 11008
rect 12176 10996 12204 11036
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 15010 11024 15016 11076
rect 15068 11024 15074 11076
rect 15212 11036 15502 11064
rect 15212 11008 15240 11036
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17405 11067 17463 11073
rect 17405 11064 17417 11067
rect 17368 11036 17417 11064
rect 17368 11024 17374 11036
rect 17405 11033 17417 11036
rect 17451 11033 17463 11067
rect 17862 11064 17868 11076
rect 17405 11027 17463 11033
rect 17512 11036 17868 11064
rect 12434 10996 12440 11008
rect 12176 10968 12440 10996
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 16761 10999 16819 11005
rect 16761 10996 16773 10999
rect 15252 10968 16773 10996
rect 15252 10956 15258 10968
rect 16761 10965 16773 10968
rect 16807 10996 16819 10999
rect 17512 10996 17540 11036
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 19760 11036 20269 11064
rect 19760 11024 19766 11036
rect 20257 11033 20269 11036
rect 20303 11064 20315 11067
rect 20916 11064 20944 11095
rect 31294 11092 31300 11144
rect 31352 11132 31358 11144
rect 31757 11135 31815 11141
rect 31757 11132 31769 11135
rect 31352 11104 31769 11132
rect 31352 11092 31358 11104
rect 31757 11101 31769 11104
rect 31803 11132 31815 11135
rect 47854 11132 47860 11144
rect 31803 11104 47860 11132
rect 31803 11101 31815 11104
rect 31757 11095 31815 11101
rect 47854 11092 47860 11104
rect 47912 11092 47918 11144
rect 20303 11036 20944 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 21726 11024 21732 11076
rect 21784 11024 21790 11076
rect 27798 11024 27804 11076
rect 27856 11064 27862 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 27856 11036 30021 11064
rect 27856 11024 27862 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 30098 11024 30104 11076
rect 30156 11064 30162 11076
rect 30156 11036 30498 11064
rect 30156 11024 30162 11036
rect 16807 10968 17540 10996
rect 16807 10965 16819 10968
rect 16761 10959 16819 10965
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 18414 10996 18420 11008
rect 17828 10968 18420 10996
rect 17828 10956 17834 10968
rect 18414 10956 18420 10968
rect 18472 10996 18478 11008
rect 20622 10996 20628 11008
rect 18472 10968 20628 10996
rect 18472 10956 18478 10968
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 3602 10792 3608 10804
rect 2148 10764 3608 10792
rect 2148 10665 2176 10764
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5859 10764 9076 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6549 10727 6607 10733
rect 6549 10693 6561 10727
rect 6595 10724 6607 10727
rect 6730 10724 6736 10736
rect 6595 10696 6736 10724
rect 6595 10693 6607 10696
rect 6549 10687 6607 10693
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 8294 10684 8300 10736
rect 8352 10684 8358 10736
rect 9048 10724 9076 10764
rect 9950 10752 9956 10804
rect 10008 10752 10014 10804
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 10962 10792 10968 10804
rect 10827 10764 10968 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 12250 10792 12256 10804
rect 11572 10764 12256 10792
rect 11572 10752 11578 10764
rect 12250 10752 12256 10764
rect 12308 10792 12314 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 12308 10764 13829 10792
rect 12308 10752 12314 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 13817 10755 13875 10761
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10761 14427 10795
rect 14369 10755 14427 10761
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15286 10792 15292 10804
rect 14875 10764 15292 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 10689 10727 10747 10733
rect 10689 10724 10701 10727
rect 9048 10696 10701 10724
rect 10689 10693 10701 10696
rect 10735 10693 10747 10727
rect 10689 10687 10747 10693
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12345 10727 12403 10733
rect 12345 10724 12357 10727
rect 12124 10696 12357 10724
rect 12124 10684 12130 10696
rect 12345 10693 12357 10696
rect 12391 10693 12403 10727
rect 14384 10724 14412 10755
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17092 10764 19257 10792
rect 17092 10752 17098 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 21450 10792 21456 10804
rect 19245 10755 19303 10761
rect 19628 10764 21456 10792
rect 15654 10724 15660 10736
rect 14384 10696 15660 10724
rect 12345 10687 12403 10693
rect 15654 10684 15660 10696
rect 15712 10684 15718 10736
rect 15746 10684 15752 10736
rect 15804 10724 15810 10736
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 15804 10696 17785 10724
rect 15804 10684 15810 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2406 10616 2412 10668
rect 2464 10616 2470 10668
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 5258 10656 5264 10668
rect 3467 10628 5264 10656
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5350 10616 5356 10668
rect 5408 10616 5414 10668
rect 7006 10616 7012 10668
rect 7064 10616 7070 10668
rect 13446 10616 13452 10668
rect 13504 10616 13510 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 4982 10588 4988 10600
rect 3743 10560 4988 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 7374 10548 7380 10600
rect 7432 10548 7438 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8110 10588 8116 10600
rect 7791 10560 8116 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7392 10520 7420 10548
rect 7064 10492 7420 10520
rect 7064 10480 7070 10492
rect 5166 10412 5172 10464
rect 5224 10412 5230 10464
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 7374 10452 7380 10464
rect 6871 10424 7380 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7484 10452 7512 10551
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 8812 10560 9505 10588
rect 8812 10548 8818 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10100 10560 10885 10588
rect 10100 10548 10106 10560
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11296 10560 12081 10588
rect 11296 10548 11302 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 14752 10588 14780 10619
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 15436 10628 15945 10656
rect 15436 10616 15442 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 12400 10560 14780 10588
rect 15013 10591 15071 10597
rect 12400 10548 12406 10560
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15194 10588 15200 10600
rect 15059 10560 15200 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 10321 10523 10379 10529
rect 10321 10520 10333 10523
rect 8772 10492 10333 10520
rect 7834 10452 7840 10464
rect 7484 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8772 10452 8800 10492
rect 10321 10489 10333 10492
rect 10367 10489 10379 10523
rect 10321 10483 10379 10489
rect 14826 10480 14832 10532
rect 14884 10520 14890 10532
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 14884 10492 15577 10520
rect 14884 10480 14890 10492
rect 15565 10489 15577 10492
rect 15611 10489 15623 10523
rect 16040 10520 16068 10551
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16356 10560 16865 10588
rect 16356 10548 16362 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 17420 10588 17448 10696
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 17773 10687 17831 10693
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 17920 10696 18262 10724
rect 17920 10684 17926 10696
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 19628 10588 19656 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21726 10752 21732 10804
rect 21784 10792 21790 10804
rect 21821 10795 21879 10801
rect 21821 10792 21833 10795
rect 21784 10764 21833 10792
rect 21784 10752 21790 10764
rect 21821 10761 21833 10764
rect 21867 10792 21879 10795
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 21867 10764 22017 10792
rect 21867 10761 21879 10764
rect 21821 10755 21879 10761
rect 22005 10761 22017 10764
rect 22051 10761 22063 10795
rect 22005 10755 22063 10761
rect 21744 10724 21772 10752
rect 21206 10696 21772 10724
rect 17420 10560 19656 10588
rect 16853 10551 16911 10557
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 22830 10588 22836 10600
rect 20027 10560 22836 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 16040 10492 16160 10520
rect 15565 10483 15623 10489
rect 8260 10424 8800 10452
rect 8260 10412 8266 10424
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 9490 10452 9496 10464
rect 9088 10424 9496 10452
rect 9088 10412 9094 10424
rect 9490 10412 9496 10424
rect 9548 10452 9554 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9548 10424 9781 10452
rect 9548 10412 9554 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 9769 10415 9827 10421
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 10560 10424 11529 10452
rect 10560 10412 10566 10424
rect 11517 10421 11529 10424
rect 11563 10452 11575 10455
rect 13998 10452 14004 10464
rect 11563 10424 14004 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 16132 10452 16160 10492
rect 20530 10452 20536 10464
rect 16132 10424 20536 10452
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 20622 10412 20628 10464
rect 20680 10452 20686 10464
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 20680 10424 21465 10452
rect 20680 10412 20686 10424
rect 21453 10421 21465 10424
rect 21499 10421 21511 10455
rect 21453 10415 21511 10421
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3786 10248 3792 10260
rect 3283 10220 3792 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 6549 10251 6607 10257
rect 6549 10217 6561 10251
rect 6595 10248 6607 10251
rect 6730 10248 6736 10260
rect 6595 10220 6736 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 6730 10208 6736 10220
rect 6788 10248 6794 10260
rect 7558 10248 7564 10260
rect 6788 10220 7564 10248
rect 6788 10208 6794 10220
rect 7558 10208 7564 10220
rect 7616 10248 7622 10260
rect 9030 10248 9036 10260
rect 7616 10220 9036 10248
rect 7616 10208 7622 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10778 10248 10784 10260
rect 10091 10220 10784 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 22278 10248 22284 10260
rect 11020 10220 22284 10248
rect 11020 10208 11026 10220
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8168 10152 8585 10180
rect 8168 10140 8174 10152
rect 8573 10149 8585 10152
rect 8619 10180 8631 10183
rect 10870 10180 10876 10192
rect 8619 10152 10876 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 13446 10140 13452 10192
rect 13504 10180 13510 10192
rect 13814 10180 13820 10192
rect 13504 10152 13820 10180
rect 13504 10140 13510 10152
rect 13814 10140 13820 10152
rect 13872 10180 13878 10192
rect 14093 10183 14151 10189
rect 14093 10180 14105 10183
rect 13872 10152 14105 10180
rect 13872 10140 13878 10152
rect 14093 10149 14105 10152
rect 14139 10149 14151 10183
rect 14093 10143 14151 10149
rect 18877 10183 18935 10189
rect 18877 10149 18889 10183
rect 18923 10180 18935 10183
rect 19150 10180 19156 10192
rect 18923 10152 19156 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 1578 10072 1584 10124
rect 1636 10072 1642 10124
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 3694 10112 3700 10124
rect 1903 10084 3700 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 3936 10084 4537 10112
rect 3936 10072 3942 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 5810 10072 5816 10124
rect 5868 10072 5874 10124
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7834 10112 7840 10124
rect 6880 10084 7840 10112
rect 6880 10072 6886 10084
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 10502 10072 10508 10124
rect 10560 10072 10566 10124
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 11974 10112 11980 10124
rect 10735 10084 11980 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3421 10047 3479 10053
rect 3421 10044 3433 10047
rect 3191 10016 3433 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3421 10013 3433 10016
rect 3467 10044 3479 10047
rect 4062 10044 4068 10056
rect 3467 10016 4068 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4430 10044 4436 10056
rect 4295 10016 4436 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4430 10004 4436 10016
rect 4488 10004 4494 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9447 10016 11100 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 3786 9936 3792 9988
rect 3844 9976 3850 9988
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 3844 9948 3985 9976
rect 3844 9936 3850 9948
rect 3973 9945 3985 9948
rect 4019 9976 4031 9979
rect 7101 9979 7159 9985
rect 4019 9948 6684 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 6656 9908 6684 9948
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7190 9976 7196 9988
rect 7147 9948 7196 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 7558 9936 7564 9988
rect 7616 9936 7622 9988
rect 10962 9976 10968 9988
rect 8404 9948 10968 9976
rect 8404 9908 8432 9948
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 6656 9880 8432 9908
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 9180 9880 10425 9908
rect 9180 9868 9186 9880
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 11072 9908 11100 10016
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 13464 10044 13492 10140
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 12650 10016 13492 10044
rect 11514 9936 11520 9988
rect 11572 9936 11578 9988
rect 14108 9976 14136 10143
rect 19150 10140 19156 10152
rect 19208 10140 19214 10192
rect 21545 10183 21603 10189
rect 21545 10149 21557 10183
rect 21591 10180 21603 10183
rect 21726 10180 21732 10192
rect 21591 10152 21732 10180
rect 21591 10149 21603 10152
rect 21545 10143 21603 10149
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 15194 10112 15200 10124
rect 14875 10084 15200 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15194 10072 15200 10084
rect 15252 10112 15258 10124
rect 16206 10112 16212 10124
rect 15252 10084 16212 10112
rect 15252 10072 15258 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17144 10084 19441 10112
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14516 10016 14565 10044
rect 14516 10004 14522 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17144 10053 17172 10084
rect 19429 10081 19441 10084
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 20162 10072 20168 10124
rect 20220 10112 20226 10124
rect 20220 10084 20852 10112
rect 20220 10072 20226 10084
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16908 10016 17141 10044
rect 16908 10004 16914 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 20824 10044 20852 10084
rect 21560 10044 21588 10143
rect 21726 10140 21732 10152
rect 21784 10140 21790 10192
rect 20824 10030 21588 10044
rect 20838 10016 21588 10030
rect 17129 10007 17187 10013
rect 15286 9976 15292 9988
rect 14108 9948 15292 9976
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 17092 9948 17417 9976
rect 17092 9936 17098 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 17512 9948 17894 9976
rect 11790 9908 11796 9920
rect 11072 9880 11796 9908
rect 10413 9871 10471 9877
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 11940 9880 13001 9908
rect 11940 9868 11946 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 16301 9911 16359 9917
rect 16301 9908 16313 9911
rect 15068 9880 16313 9908
rect 15068 9868 15074 9880
rect 16301 9877 16313 9880
rect 16347 9877 16359 9911
rect 16301 9871 16359 9877
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16577 9911 16635 9917
rect 16577 9908 16589 9911
rect 16540 9880 16589 9908
rect 16540 9868 16546 9880
rect 16577 9877 16589 9880
rect 16623 9908 16635 9911
rect 16761 9911 16819 9917
rect 16761 9908 16773 9911
rect 16623 9880 16773 9908
rect 16623 9877 16635 9880
rect 16577 9871 16635 9877
rect 16761 9877 16773 9880
rect 16807 9908 16819 9911
rect 17512 9908 17540 9948
rect 16807 9880 17540 9908
rect 17788 9908 17816 9948
rect 19702 9936 19708 9988
rect 19760 9936 19766 9988
rect 24118 9976 24124 9988
rect 21008 9948 24124 9976
rect 18322 9908 18328 9920
rect 17788 9880 18328 9908
rect 16807 9877 16819 9880
rect 16761 9871 16819 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 19720 9908 19748 9936
rect 21008 9908 21036 9948
rect 24118 9936 24124 9948
rect 24176 9936 24182 9988
rect 19720 9880 21036 9908
rect 21174 9868 21180 9920
rect 21232 9868 21238 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1486 9664 1492 9716
rect 1544 9664 1550 9716
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 13630 9704 13636 9716
rect 7432 9676 13636 9704
rect 7432 9664 7438 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 13814 9704 13820 9716
rect 13740 9676 13820 9704
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5767 9608 5825 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 5813 9605 5825 9608
rect 5859 9636 5871 9639
rect 5994 9636 6000 9648
rect 5859 9608 6000 9636
rect 5859 9605 5871 9608
rect 5813 9599 5871 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 8389 9639 8447 9645
rect 8389 9605 8401 9639
rect 8435 9636 8447 9639
rect 8662 9636 8668 9648
rect 8435 9608 8668 9636
rect 8435 9605 8447 9608
rect 8389 9599 8447 9605
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 13740 9636 13768 9676
rect 13814 9664 13820 9676
rect 13872 9704 13878 9716
rect 13909 9707 13967 9713
rect 13909 9704 13921 9707
rect 13872 9676 13921 9704
rect 13872 9664 13878 9676
rect 13909 9673 13921 9676
rect 13955 9673 13967 9707
rect 13909 9667 13967 9673
rect 16206 9664 16212 9716
rect 16264 9664 16270 9716
rect 18414 9704 18420 9716
rect 17512 9676 18420 9704
rect 16482 9636 16488 9648
rect 13202 9608 13768 9636
rect 15962 9608 16488 9636
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17512 9636 17540 9676
rect 18414 9664 18420 9676
rect 18472 9704 18478 9716
rect 19150 9704 19156 9716
rect 18472 9676 19156 9704
rect 18472 9664 18478 9676
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 18690 9636 18696 9648
rect 17175 9608 17540 9636
rect 18354 9608 18696 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 18690 9596 18696 9608
rect 18748 9596 18754 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 24578 9636 24584 9648
rect 19567 9608 24584 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 24578 9596 24584 9608
rect 24636 9596 24642 9648
rect 28445 9639 28503 9645
rect 28445 9605 28457 9639
rect 28491 9636 28503 9639
rect 31294 9636 31300 9648
rect 28491 9608 31300 9636
rect 28491 9605 28503 9608
rect 28445 9599 28503 9605
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 3786 9528 3792 9580
rect 3844 9528 3850 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 5166 9568 5172 9580
rect 4295 9540 5172 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8120 9572 8178 9577
rect 8036 9571 8178 9572
rect 8036 9568 8132 9571
rect 7892 9544 8132 9568
rect 7892 9540 8064 9544
rect 7892 9528 7898 9540
rect 8120 9537 8132 9544
rect 8166 9537 8178 9571
rect 8120 9531 8178 9537
rect 9490 9528 9496 9580
rect 9548 9528 9554 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9732 9540 10701 9568
rect 9732 9528 9738 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1728 9472 1961 9500
rect 1728 9460 1734 9472
rect 1949 9469 1961 9472
rect 1995 9500 2007 9503
rect 2590 9500 2596 9512
rect 1995 9472 2596 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 4522 9460 4528 9512
rect 4580 9460 4586 9512
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 6822 9500 6828 9512
rect 6779 9472 6828 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7742 9460 7748 9512
rect 7800 9500 7806 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 7800 9472 10793 9500
rect 7800 9460 7806 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11296 9472 11713 9500
rect 11296 9460 11302 9472
rect 11701 9469 11713 9472
rect 11747 9500 11759 9503
rect 14458 9500 14464 9512
rect 11747 9472 14464 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 14568 9472 14749 9500
rect 3602 9392 3608 9444
rect 3660 9392 3666 9444
rect 13538 9392 13544 9444
rect 13596 9432 13602 9444
rect 14568 9432 14596 9472
rect 14737 9469 14749 9472
rect 14783 9500 14795 9503
rect 16666 9500 16672 9512
rect 14783 9472 16672 9500
rect 14783 9469 14795 9472
rect 14737 9463 14795 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17126 9500 17132 9512
rect 16960 9472 17132 9500
rect 16960 9432 16988 9472
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 19444 9500 19472 9531
rect 27522 9528 27528 9580
rect 27580 9528 27586 9580
rect 17276 9472 19472 9500
rect 19705 9503 19763 9509
rect 17276 9460 17282 9472
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21174 9500 21180 9512
rect 19751 9472 21180 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 22612 9472 27997 9500
rect 22612 9460 22618 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 13596 9404 14596 9432
rect 16040 9404 16988 9432
rect 13596 9392 13602 9404
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 8754 9364 8760 9376
rect 7248 9336 8760 9364
rect 7248 9324 7254 9336
rect 8754 9324 8760 9336
rect 8812 9364 8818 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8812 9336 9873 9364
rect 8812 9324 8818 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 11606 9364 11612 9376
rect 10367 9336 11612 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 12492 9336 13461 9364
rect 12492 9324 12498 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 16040 9364 16068 9404
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 18380 9404 18736 9432
rect 18380 9392 18386 9404
rect 18708 9376 18736 9404
rect 19058 9392 19064 9444
rect 19116 9392 19122 9444
rect 14608 9336 16068 9364
rect 14608 9324 14614 9336
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 16172 9336 18613 9364
rect 16172 9324 16178 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18601 9327 18659 9333
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 18748 9336 20085 9364
rect 18748 9324 18754 9336
rect 20073 9333 20085 9336
rect 20119 9364 20131 9367
rect 20162 9364 20168 9376
rect 20119 9336 20168 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 27801 9367 27859 9373
rect 27801 9333 27813 9367
rect 27847 9364 27859 9367
rect 28460 9364 28488 9599
rect 31294 9596 31300 9608
rect 31352 9596 31358 9648
rect 27847 9336 28488 9364
rect 27847 9333 27859 9336
rect 27801 9327 27859 9333
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 2740 9132 3801 9160
rect 2740 9120 2746 9132
rect 3789 9129 3801 9132
rect 3835 9160 3847 9163
rect 3835 9132 4016 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 1578 8984 1584 9036
rect 1636 8984 1642 9036
rect 3988 9033 4016 9132
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 4672 9132 4752 9160
rect 4672 9120 4678 9132
rect 4724 9033 4752 9132
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 9674 9160 9680 9172
rect 7883 9132 9680 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10134 9120 10140 9172
rect 10192 9120 10198 9172
rect 11563 9163 11621 9169
rect 11563 9129 11575 9163
rect 11609 9160 11621 9163
rect 32858 9160 32864 9172
rect 11609 9132 32864 9160
rect 11609 9129 11621 9132
rect 11563 9123 11621 9129
rect 32858 9120 32864 9132
rect 32916 9120 32922 9172
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 6880 9064 8340 9092
rect 6880 9052 6886 9064
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 3973 9027 4031 9033
rect 1903 8996 3924 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2924 8928 3065 8956
rect 2924 8916 2930 8928
rect 3053 8925 3065 8928
rect 3099 8956 3111 8959
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3099 8928 3341 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3896 8956 3924 8996
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 5534 8956 5540 8968
rect 3896 8928 5540 8956
rect 3329 8919 3387 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7742 8956 7748 8968
rect 7423 8928 7748 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 5920 8888 5948 8919
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 7984 8928 8217 8956
rect 7984 8916 7990 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8312 8956 8340 9064
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 10042 9092 10048 9104
rect 8720 9064 10048 9092
rect 8720 9052 8726 9064
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 11974 9092 11980 9104
rect 10704 9064 11980 9092
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 9024 8447 9027
rect 8754 9024 8760 9036
rect 8435 8996 8760 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 10704 9024 10732 9064
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 14277 9095 14335 9101
rect 14277 9061 14289 9095
rect 14323 9092 14335 9095
rect 14734 9092 14740 9104
rect 14323 9064 14740 9092
rect 14323 9061 14335 9064
rect 14277 9055 14335 9061
rect 14734 9052 14740 9064
rect 14792 9052 14798 9104
rect 15470 9092 15476 9104
rect 14844 9064 15476 9092
rect 9640 8996 10732 9024
rect 10781 9027 10839 9033
rect 9640 8984 9646 8996
rect 10781 8993 10793 9027
rect 10827 9024 10839 9027
rect 10827 8996 11744 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 10226 8956 10232 8968
rect 8312 8928 10232 8956
rect 8205 8919 8263 8925
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10376 8928 11345 8956
rect 10376 8916 10382 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11716 8956 11744 8996
rect 11790 8984 11796 9036
rect 11848 9024 11854 9036
rect 14844 9024 14872 9064
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 11848 8996 14872 9024
rect 14921 9027 14979 9033
rect 11848 8984 11854 8996
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15746 9024 15752 9036
rect 14967 8996 15752 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 11716 8928 13308 8956
rect 11333 8919 11391 8925
rect 9122 8888 9128 8900
rect 5920 8860 9128 8888
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 9490 8888 9496 8900
rect 9232 8860 9496 8888
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 6638 8820 6644 8832
rect 2915 8792 6644 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9232 8820 9260 8860
rect 9490 8848 9496 8860
rect 9548 8888 9554 8900
rect 10042 8888 10048 8900
rect 9548 8860 10048 8888
rect 9548 8848 9554 8860
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 10505 8891 10563 8897
rect 10505 8857 10517 8891
rect 10551 8888 10563 8891
rect 11882 8888 11888 8900
rect 10551 8860 11888 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 13170 8888 13176 8900
rect 12032 8860 13176 8888
rect 12032 8848 12038 8860
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 9079 8792 9260 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 9732 8792 10609 8820
rect 9732 8780 9738 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12584 8792 12633 8820
rect 12584 8780 12590 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 13280 8820 13308 8928
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 14737 8959 14795 8965
rect 14737 8956 14749 8959
rect 13412 8928 14749 8956
rect 13412 8916 13418 8928
rect 14737 8925 14749 8928
rect 14783 8925 14795 8959
rect 14737 8919 14795 8925
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 13587 8860 14657 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 14645 8851 14703 8857
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 16264 8860 16313 8888
rect 16264 8848 16270 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 17526 8860 18184 8888
rect 16301 8851 16359 8857
rect 15010 8820 15016 8832
rect 13280 8792 15016 8820
rect 12621 8783 12679 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17586 8820 17592 8832
rect 16724 8792 17592 8820
rect 16724 8780 16730 8792
rect 17586 8780 17592 8792
rect 17644 8820 17650 8832
rect 18156 8829 18184 8860
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17644 8792 17785 8820
rect 17644 8780 17650 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18690 8820 18696 8832
rect 18187 8792 18696 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18690 8780 18696 8792
rect 18748 8820 18754 8832
rect 18969 8823 19027 8829
rect 18969 8820 18981 8823
rect 18748 8792 18981 8820
rect 18748 8780 18754 8792
rect 18969 8789 18981 8792
rect 19015 8789 19027 8823
rect 18969 8783 19027 8789
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 3326 8576 3332 8628
rect 3384 8576 3390 8628
rect 3970 8576 3976 8628
rect 4028 8576 4034 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5316 8588 5825 8616
rect 5316 8576 5322 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 7282 8576 7288 8628
rect 7340 8576 7346 8628
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 9582 8616 9588 8628
rect 7432 8588 9588 8616
rect 7432 8576 7438 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 12342 8616 12348 8628
rect 10183 8588 12348 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12526 8576 12532 8628
rect 12584 8576 12590 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 15378 8616 15384 8628
rect 14323 8588 15384 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8585 15623 8619
rect 15565 8579 15623 8585
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16298 8616 16304 8628
rect 15979 8588 16304 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 3513 8551 3571 8557
rect 3513 8548 3525 8551
rect 2792 8520 3525 8548
rect 2792 8492 2820 8520
rect 3513 8517 3525 8520
rect 3559 8517 3571 8551
rect 3513 8511 3571 8517
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 5350 8548 5356 8560
rect 5224 8520 5356 8548
rect 5224 8508 5230 8520
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 7193 8551 7251 8557
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 11790 8548 11796 8560
rect 7239 8520 11796 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 15580 8548 15608 8579
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 20438 8548 20444 8560
rect 15580 8520 20444 8548
rect 20438 8508 20444 8520
rect 20496 8508 20502 8560
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 2774 8480 2780 8492
rect 1627 8452 2780 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3326 8480 3332 8492
rect 3099 8452 3332 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 4982 8480 4988 8492
rect 4847 8452 4988 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 6362 8480 6368 8492
rect 6043 8452 6368 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 8312 8452 8524 8480
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 6454 8412 6460 8424
rect 1903 8384 6460 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 8312 8412 8340 8452
rect 6840 8384 8340 8412
rect 8389 8415 8447 8421
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 4338 8344 4344 8356
rect 2915 8316 4344 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 6840 8344 6868 8384
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8496 8412 8524 8452
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8628 8452 8677 8480
rect 8628 8440 8634 8452
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 13538 8480 13544 8492
rect 10796 8452 13544 8480
rect 8496 8384 9720 8412
rect 8389 8375 8447 8381
rect 4663 8316 6868 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 8404 8344 8432 8375
rect 9582 8344 9588 8356
rect 6972 8316 8340 8344
rect 8404 8316 9588 8344
rect 6972 8304 6978 8316
rect 8312 8276 8340 8316
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 9692 8344 9720 8384
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 10796 8421 10824 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13679 8452 14657 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 18414 8480 18420 8492
rect 14645 8443 14703 8449
rect 14936 8452 18420 8480
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 14550 8412 14556 8424
rect 12851 8384 14556 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14734 8372 14740 8424
rect 14792 8372 14798 8424
rect 14936 8421 14964 8452
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 20346 8412 20352 8424
rect 16255 8384 20352 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 11054 8344 11060 8356
rect 9692 8316 11060 8344
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 12161 8347 12219 8353
rect 11164 8316 12112 8344
rect 11164 8276 11192 8316
rect 8312 8248 11192 8276
rect 12084 8276 12112 8316
rect 12161 8313 12173 8347
rect 12207 8344 12219 8347
rect 12434 8344 12440 8356
rect 12207 8316 12440 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 16040 8344 16068 8375
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 12544 8316 16068 8344
rect 12544 8276 12572 8316
rect 12084 8248 12572 8276
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 14734 8276 14740 8288
rect 13412 8248 14740 8276
rect 13412 8236 13418 8248
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1670 8072 1676 8084
rect 1627 8044 1676 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3476 8044 3801 8072
rect 3476 8032 3482 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4212 8044 4353 8072
rect 4212 8032 4218 8044
rect 4341 8041 4353 8044
rect 4387 8072 4399 8075
rect 4387 8044 7144 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 7116 8004 7144 8044
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 8352 8044 9597 8072
rect 8352 8032 8358 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 12989 8075 13047 8081
rect 10008 8044 11836 8072
rect 10008 8032 10014 8044
rect 8386 8004 8392 8016
rect 2915 7976 7052 8004
rect 7116 7976 8392 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 2746 7908 3525 7936
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2746 7868 2774 7908
rect 3513 7905 3525 7908
rect 3559 7936 3571 7939
rect 3694 7936 3700 7948
rect 3559 7908 3700 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 2455 7840 2774 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 1780 7800 1808 7831
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2924 7840 3065 7868
rect 2924 7828 2930 7840
rect 3053 7837 3065 7840
rect 3099 7868 3111 7871
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3099 7840 3341 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 7024 7868 7052 7976
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 11698 8004 11704 8016
rect 10060 7976 11704 8004
rect 10060 7945 10088 7976
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 10134 7896 10140 7948
rect 10192 7896 10198 7948
rect 11146 7896 11152 7948
rect 11204 7896 11210 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 11388 7908 11529 7936
rect 11388 7896 11394 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11808 7936 11836 8044
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 17218 8072 17224 8084
rect 13035 8044 17224 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12032 7976 15056 8004
rect 12032 7964 12038 7976
rect 13354 7936 13360 7948
rect 11808 7908 13360 7936
rect 11517 7899 11575 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 13587 7908 13676 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 11164 7868 11192 7896
rect 7024 7840 11192 7868
rect 11241 7871 11299 7877
rect 3329 7831 3387 7837
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 3418 7800 3424 7812
rect 1780 7772 3424 7800
rect 3418 7760 3424 7772
rect 3476 7760 3482 7812
rect 11149 7803 11207 7809
rect 11149 7769 11161 7803
rect 11195 7800 11207 7803
rect 11256 7800 11284 7831
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 11480 7840 13461 7868
rect 11480 7828 11486 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 13648 7800 13676 7908
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 13780 7908 14841 7936
rect 13780 7896 13786 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15028 7877 15056 7976
rect 15194 7964 15200 8016
rect 15252 7964 15258 8016
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 22554 7868 22560 7880
rect 15059 7840 22560 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 19702 7800 19708 7812
rect 11195 7772 13492 7800
rect 13648 7772 19708 7800
rect 11195 7769 11207 7772
rect 11149 7763 11207 7769
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 6086 7732 6092 7744
rect 2271 7704 6092 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 9950 7692 9956 7744
rect 10008 7692 10014 7744
rect 13354 7692 13360 7744
rect 13412 7692 13418 7744
rect 13464 7732 13492 7772
rect 19702 7760 19708 7772
rect 19760 7760 19766 7812
rect 16574 7732 16580 7744
rect 13464 7704 16580 7732
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1946 7528 1952 7540
rect 1627 7500 1952 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 2096 7500 2237 7528
rect 2096 7488 2102 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 3326 7528 3332 7540
rect 2225 7491 2283 7497
rect 2332 7500 3332 7528
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 1854 7392 1860 7404
rect 1811 7364 1860 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 1854 7352 1860 7364
rect 1912 7392 1918 7404
rect 2332 7392 2360 7500
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 3510 7488 3516 7540
rect 3568 7488 3574 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13412 7500 13461 7528
rect 13412 7488 13418 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 27798 7528 27804 7540
rect 23992 7500 27804 7528
rect 23992 7488 23998 7500
rect 27798 7488 27804 7500
rect 27856 7488 27862 7540
rect 4157 7463 4215 7469
rect 4157 7460 4169 7463
rect 2516 7432 4169 7460
rect 2516 7404 2544 7432
rect 4157 7429 4169 7432
rect 4203 7429 4215 7463
rect 4157 7423 4215 7429
rect 9214 7420 9220 7472
rect 9272 7460 9278 7472
rect 9272 7432 10916 7460
rect 9272 7420 9278 7432
rect 1912 7364 2360 7392
rect 2409 7395 2467 7401
rect 1912 7352 1918 7364
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2498 7392 2504 7404
rect 2455 7364 2504 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7361 3111 7395
rect 3053 7355 3111 7361
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 3068 7324 3096 7355
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3752 7364 3985 7392
rect 3752 7352 3758 7364
rect 3973 7361 3985 7364
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10888 7392 10916 7432
rect 11606 7420 11612 7472
rect 11664 7460 11670 7472
rect 24026 7460 24032 7472
rect 11664 7432 14320 7460
rect 23690 7432 24032 7460
rect 11664 7420 11670 7432
rect 14292 7401 14320 7432
rect 24026 7420 24032 7432
rect 24084 7460 24090 7472
rect 24213 7463 24271 7469
rect 24213 7460 24225 7463
rect 24084 7432 24225 7460
rect 24084 7420 24090 7432
rect 24213 7429 24225 7432
rect 24259 7429 24271 7463
rect 24213 7423 24271 7429
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 10888 7364 12725 7392
rect 10781 7355 10839 7361
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 2832 7296 3096 7324
rect 2832 7284 2838 7296
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 3384 7296 4353 7324
rect 3384 7284 3390 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 10796 7324 10824 7355
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 7708 7296 10824 7324
rect 7708 7284 7714 7296
rect 22462 7284 22468 7336
rect 22520 7284 22526 7336
rect 10597 7259 10655 7265
rect 10597 7225 10609 7259
rect 10643 7256 10655 7259
rect 15654 7256 15660 7268
rect 10643 7228 15660 7256
rect 10643 7225 10655 7228
rect 10597 7219 10655 7225
rect 15654 7216 15660 7228
rect 15712 7216 15718 7268
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 9030 7188 9036 7200
rect 2915 7160 9036 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7188 12587 7191
rect 13998 7188 14004 7200
rect 12575 7160 14004 7188
rect 12575 7157 12587 7160
rect 12529 7151 12587 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 17494 7188 17500 7200
rect 14139 7160 17500 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 2225 6987 2283 6993
rect 2225 6953 2237 6987
rect 2271 6984 2283 6987
rect 23201 6987 23259 6993
rect 2271 6956 3924 6984
rect 2271 6953 2283 6956
rect 2225 6947 2283 6953
rect 2774 6876 2780 6928
rect 2832 6916 2838 6928
rect 3329 6919 3387 6925
rect 3329 6916 3341 6919
rect 2832 6888 3341 6916
rect 2832 6876 2838 6888
rect 3329 6885 3341 6888
rect 3375 6885 3387 6919
rect 3329 6879 3387 6885
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 2424 6820 3801 6848
rect 2424 6792 2452 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3896 6848 3924 6956
rect 23201 6953 23213 6987
rect 23247 6984 23259 6987
rect 23934 6984 23940 6996
rect 23247 6956 23940 6984
rect 23247 6953 23259 6956
rect 23201 6947 23259 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 8846 6848 8852 6860
rect 3896 6820 8852 6848
rect 3789 6811 3847 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2406 6740 2412 6792
rect 2464 6740 2470 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2746 6752 3065 6780
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 2746 6712 2774 6752
rect 3053 6749 3065 6752
rect 3099 6780 3111 6783
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3099 6752 3525 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 20956 6752 22937 6780
rect 20956 6740 20962 6752
rect 22925 6749 22937 6752
rect 22971 6780 22983 6783
rect 27522 6780 27528 6792
rect 22971 6752 27528 6780
rect 22971 6749 22983 6752
rect 22925 6743 22983 6749
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 10686 6712 10692 6724
rect 1360 6684 2774 6712
rect 2884 6684 10692 6712
rect 1360 6672 1366 6684
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 2884 6653 2912 6684
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1452 6616 1593 6644
rect 1452 6604 1458 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 23385 6647 23443 6653
rect 23385 6644 23397 6647
rect 22152 6616 23397 6644
rect 22152 6604 22158 6616
rect 23385 6613 23397 6616
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 3970 6440 3976 6452
rect 1820 6412 3976 6440
rect 1820 6400 1826 6412
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2924 6276 3065 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6276
rect 3099 6304 3111 6307
rect 3329 6307 3387 6313
rect 3329 6304 3341 6307
rect 3099 6276 3341 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3329 6273 3341 6276
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 22440 6307 22498 6313
rect 22440 6273 22452 6307
rect 22486 6304 22498 6307
rect 22554 6304 22560 6316
rect 22486 6276 22560 6304
rect 22486 6273 22498 6276
rect 22440 6267 22498 6273
rect 22554 6264 22560 6276
rect 22612 6264 22618 6316
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 1360 6208 1593 6236
rect 1360 6196 1366 6208
rect 1581 6205 1593 6208
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 12158 6236 12164 6248
rect 1903 6208 12164 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 7466 6168 7472 6180
rect 2915 6140 7472 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 22511 6103 22569 6109
rect 22511 6069 22523 6103
rect 22557 6100 22569 6103
rect 24854 6100 24860 6112
rect 22557 6072 24860 6100
rect 22557 6069 22569 6072
rect 22511 6063 22569 6069
rect 24854 6060 24860 6072
rect 24912 6060 24918 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 1360 5868 2697 5896
rect 1360 5856 1366 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 18923 5868 21005 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 22462 5896 22468 5908
rect 21039 5868 22468 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 12860 5800 17264 5828
rect 12860 5788 12866 5800
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 15764 5769 15792 5800
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 14056 5732 15577 5760
rect 14056 5720 14062 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16908 5732 17141 5760
rect 16908 5720 16914 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17236 5760 17264 5800
rect 22094 5760 22100 5772
rect 17236 5732 22100 5760
rect 17129 5723 17187 5729
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 24854 5720 24860 5772
rect 24912 5720 24918 5772
rect 26973 5763 27031 5769
rect 26973 5729 26985 5763
rect 27019 5760 27031 5763
rect 28718 5760 28724 5772
rect 27019 5732 28724 5760
rect 27019 5729 27031 5732
rect 26973 5723 27031 5729
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 9766 5692 9772 5704
rect 1903 5664 9772 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 1596 5624 1624 5655
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 20898 5652 20904 5704
rect 20956 5652 20962 5704
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 2869 5627 2927 5633
rect 2869 5624 2881 5627
rect 1596 5596 2881 5624
rect 2869 5593 2881 5596
rect 2915 5593 2927 5627
rect 2869 5587 2927 5593
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 16632 5596 17417 5624
rect 16632 5584 16638 5596
rect 17405 5593 17417 5596
rect 17451 5593 17463 5627
rect 18690 5624 18696 5636
rect 18630 5596 18696 5624
rect 17405 5587 17463 5593
rect 18690 5584 18696 5596
rect 18748 5624 18754 5636
rect 19337 5627 19395 5633
rect 19337 5624 19349 5627
rect 18748 5596 19349 5624
rect 18748 5584 18754 5596
rect 19337 5593 19349 5596
rect 19383 5593 19395 5627
rect 24688 5624 24716 5655
rect 25498 5624 25504 5636
rect 24688 5596 25504 5624
rect 19337 5587 19395 5593
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 26513 5627 26571 5633
rect 26513 5593 26525 5627
rect 26559 5593 26571 5627
rect 26513 5587 26571 5593
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 17034 5556 17040 5568
rect 16255 5528 17040 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 21358 5516 21364 5568
rect 21416 5516 21422 5568
rect 26528 5556 26556 5587
rect 27154 5584 27160 5636
rect 27212 5584 27218 5636
rect 27338 5584 27344 5636
rect 27396 5624 27402 5636
rect 27522 5624 27528 5636
rect 27396 5596 27528 5624
rect 27396 5584 27402 5596
rect 27522 5584 27528 5596
rect 27580 5584 27586 5636
rect 28813 5627 28871 5633
rect 28813 5593 28825 5627
rect 28859 5624 28871 5627
rect 28902 5624 28908 5636
rect 28859 5596 28908 5624
rect 28859 5593 28871 5596
rect 28813 5587 28871 5593
rect 28902 5584 28908 5596
rect 28960 5584 28966 5636
rect 27614 5556 27620 5568
rect 26528 5528 27620 5556
rect 27614 5516 27620 5528
rect 27672 5556 27678 5568
rect 28534 5556 28540 5568
rect 27672 5528 28540 5556
rect 27672 5516 27678 5528
rect 28534 5516 28540 5528
rect 28592 5516 28598 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 22879 5355 22937 5361
rect 22879 5321 22891 5355
rect 22925 5352 22937 5355
rect 27154 5352 27160 5364
rect 22925 5324 27160 5352
rect 22925 5321 22937 5324
rect 22879 5315 22937 5321
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 28350 5244 28356 5296
rect 28408 5284 28414 5296
rect 28408 5256 30328 5284
rect 28408 5244 28414 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1360 5188 1593 5216
rect 1360 5176 1366 5188
rect 1581 5185 1593 5188
rect 1627 5216 1639 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 1627 5188 2697 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 21358 5216 21364 5228
rect 17604 5188 21364 5216
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 9858 5148 9864 5160
rect 1903 5120 9864 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15528 5120 15853 5148
rect 15528 5108 15534 5120
rect 15841 5117 15853 5120
rect 15887 5148 15899 5151
rect 17604 5148 17632 5188
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 22094 5176 22100 5228
rect 22152 5225 22158 5228
rect 22152 5219 22190 5225
rect 22178 5185 22190 5219
rect 22776 5219 22834 5225
rect 22776 5216 22788 5219
rect 22152 5179 22190 5185
rect 22296 5188 22788 5216
rect 22152 5176 22158 5179
rect 15887 5120 17632 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 17678 5108 17684 5160
rect 17736 5108 17742 5160
rect 21376 5148 21404 5176
rect 22296 5148 22324 5188
rect 22776 5185 22788 5188
rect 22822 5185 22834 5219
rect 22776 5179 22834 5185
rect 21376 5120 22324 5148
rect 28629 5151 28687 5157
rect 28629 5117 28641 5151
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 28644 5080 28672 5111
rect 28810 5108 28816 5160
rect 28868 5108 28874 5160
rect 30300 5157 30328 5256
rect 30285 5151 30343 5157
rect 30285 5117 30297 5151
rect 30331 5148 30343 5151
rect 41414 5148 41420 5160
rect 30331 5120 41420 5148
rect 30331 5117 30343 5120
rect 30285 5111 30343 5117
rect 41414 5108 41420 5120
rect 41472 5108 41478 5160
rect 33502 5080 33508 5092
rect 28644 5052 33508 5080
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 17862 5012 17868 5024
rect 16347 4984 17868 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 20530 5012 20536 5024
rect 18187 4984 20536 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22235 5015 22293 5021
rect 22235 4981 22247 5015
rect 22281 5012 22293 5015
rect 25958 5012 25964 5024
rect 22281 4984 25964 5012
rect 22281 4981 22293 4984
rect 22235 4975 22293 4981
rect 25958 4972 25964 4984
rect 26016 4972 26022 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 16632 4780 19533 4808
rect 16632 4768 16638 4780
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 24719 4811 24777 4817
rect 24719 4777 24731 4811
rect 24765 4808 24777 4811
rect 28810 4808 28816 4820
rect 24765 4780 28816 4808
rect 24765 4777 24777 4780
rect 24719 4771 24777 4777
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 1360 4644 1593 4672
rect 1360 4632 1366 4644
rect 1581 4641 1593 4644
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 11514 4672 11520 4684
rect 1903 4644 11520 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1596 4604 1624 4635
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 25958 4632 25964 4684
rect 26016 4632 26022 4684
rect 27522 4632 27528 4684
rect 27580 4632 27586 4684
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 1596 4576 2881 4604
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20898 4604 20904 4616
rect 19475 4576 20904 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 22066 4576 24628 4604
rect 2774 4428 2780 4480
rect 2832 4428 2838 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 17736 4440 19901 4468
rect 17736 4428 17742 4440
rect 19889 4437 19901 4440
rect 19935 4468 19947 4471
rect 22066 4468 22094 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 25777 4607 25835 4613
rect 25777 4573 25789 4607
rect 25823 4573 25835 4607
rect 25777 4567 25835 4573
rect 19935 4440 22094 4468
rect 25792 4468 25820 4567
rect 27798 4468 27804 4480
rect 25792 4440 27804 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 27798 4428 27804 4440
rect 27856 4428 27862 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2271 4236 2912 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2774 4156 2780 4208
rect 2832 4156 2838 4208
rect 2884 4196 2912 4236
rect 2884 4168 3464 4196
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2792 4128 2820 4156
rect 2455 4100 2820 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2924 4100 3065 4128
rect 2924 4088 2930 4100
rect 3053 4097 3065 4100
rect 3099 4128 3111 4131
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3099 4100 3341 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 2869 3995 2927 4001
rect 2869 3992 2881 3995
rect 2740 3964 2881 3992
rect 2740 3952 2746 3964
rect 2869 3961 2881 3964
rect 2915 3961 2927 3995
rect 3436 3992 3464 4168
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 10594 4128 10600 4140
rect 6328 4100 10600 4128
rect 6328 4088 6334 4100
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 9950 3992 9956 4004
rect 3436 3964 9956 3992
rect 2869 3955 2927 3961
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 9674 3924 9680 3936
rect 1627 3896 9680 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 1302 3680 1308 3732
rect 1360 3720 1366 3732
rect 2774 3720 2780 3732
rect 1360 3692 2780 3720
rect 1360 3680 1366 3692
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 11422 3720 11428 3732
rect 2915 3692 11428 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 3513 3655 3571 3661
rect 3513 3652 3525 3655
rect 2608 3624 3525 3652
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3516 1639 3519
rect 2608 3516 2636 3624
rect 3513 3621 3525 3624
rect 3559 3621 3571 3655
rect 3513 3615 3571 3621
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 44082 3652 44088 3664
rect 28960 3624 44088 3652
rect 28960 3612 28966 3624
rect 44082 3612 44088 3624
rect 44140 3612 44146 3664
rect 7006 3584 7012 3596
rect 1627 3488 2636 3516
rect 2746 3556 7012 3584
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1811 3383 1869 3389
rect 1811 3349 1823 3383
rect 1857 3380 1869 3383
rect 2746 3380 2774 3556
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 27522 3544 27528 3596
rect 27580 3584 27586 3596
rect 46750 3584 46756 3596
rect 27580 3556 46756 3584
rect 27580 3544 27586 3556
rect 46750 3544 46756 3556
rect 46808 3544 46814 3596
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 11517 3519 11575 3525
rect 3099 3488 3372 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3344 3392 3372 3488
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11974 3516 11980 3528
rect 11563 3488 11980 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 28534 3476 28540 3528
rect 28592 3516 28598 3528
rect 49418 3516 49424 3528
rect 28592 3488 49424 3516
rect 28592 3476 28598 3488
rect 49418 3476 49424 3488
rect 49476 3476 49482 3528
rect 3418 3408 3424 3460
rect 3476 3448 3482 3460
rect 12618 3448 12624 3460
rect 3476 3420 12624 3448
rect 3476 3408 3482 3420
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 38746 3448 38752 3460
rect 19392 3420 38752 3448
rect 19392 3408 19398 3420
rect 38746 3408 38752 3420
rect 38804 3408 38810 3460
rect 1857 3352 2774 3380
rect 1857 3349 1869 3352
rect 1811 3343 1869 3349
rect 3326 3340 3332 3392
rect 3384 3340 3390 3392
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3418 3176 3424 3188
rect 2915 3148 3424 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 8352 3148 12725 3176
rect 8352 3136 8358 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 12713 3139 12771 3145
rect 6914 3108 6920 3120
rect 1872 3080 6920 3108
rect 1872 3049 1900 3080
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 10042 3068 10048 3120
rect 10100 3068 10106 3120
rect 12621 3111 12679 3117
rect 12621 3077 12633 3111
rect 12667 3108 12679 3111
rect 12802 3108 12808 3120
rect 12667 3080 12808 3108
rect 12667 3077 12679 3080
rect 12621 3071 12679 3077
rect 12802 3068 12808 3080
rect 12860 3068 12866 3120
rect 13909 3111 13967 3117
rect 13909 3077 13921 3111
rect 13955 3108 13967 3111
rect 15470 3108 15476 3120
rect 13955 3080 15476 3108
rect 13955 3077 13967 3080
rect 13909 3071 13967 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 17678 3108 17684 3120
rect 15611 3080 17684 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2832 3012 3065 3040
rect 2832 3000 2838 3012
rect 3053 3009 3065 3012
rect 3099 3040 3111 3043
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 3099 3012 3341 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7892 3012 8769 3040
rect 7892 3000 7898 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17920 3012 18337 3040
rect 17920 3000 17926 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20530 3000 20536 3052
rect 20588 3000 20594 3052
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1360 2944 1593 2972
rect 1360 2932 1366 2944
rect 1581 2941 1593 2944
rect 1627 2972 1639 2975
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 1627 2944 3525 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 7248 2944 9045 2972
rect 7248 2932 7254 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 9824 2944 14105 2972
rect 9824 2932 9830 2944
rect 14093 2941 14105 2944
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 10551 2876 11468 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 2866 2836 2872 2848
rect 1452 2808 2872 2836
rect 1452 2796 1458 2808
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 10100 2808 10793 2836
rect 10100 2796 10106 2808
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 11440 2836 11468 2876
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 12492 2876 15761 2904
rect 12492 2864 12498 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 16574 2836 16580 2848
rect 11440 2808 16580 2836
rect 10781 2799 10839 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17494 2836 17500 2848
rect 16899 2808 17500 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 20070 2836 20076 2848
rect 18187 2808 20076 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20349 2839 20407 2845
rect 20349 2805 20361 2839
rect 20395 2836 20407 2839
rect 22002 2836 22008 2848
rect 20395 2808 22008 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 7190 2632 7196 2644
rect 2915 2604 7196 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27856 2604 28181 2632
rect 27856 2592 27862 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 28776 2604 30849 2632
rect 28776 2592 28782 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 33502 2592 33508 2644
rect 33560 2592 33566 2644
rect 11606 2564 11612 2576
rect 5552 2536 11612 2564
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1360 2468 1593 2496
rect 1360 2456 1366 2468
rect 1581 2465 1593 2468
rect 1627 2496 1639 2499
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 1627 2468 3525 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 3513 2465 3525 2468
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 1872 2360 1900 2391
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2924 2400 3065 2428
rect 2924 2388 2930 2400
rect 3053 2397 3065 2400
rect 3099 2428 3111 2431
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3099 2400 3341 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 5552 2428 5580 2536
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 14792 2468 15301 2496
rect 14792 2456 14798 2468
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17460 2468 17969 2496
rect 17460 2456 17466 2468
rect 17957 2465 17969 2468
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22796 2468 23121 2496
rect 22796 2456 22802 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 27338 2456 27344 2508
rect 27396 2496 27402 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 27396 2468 36369 2496
rect 27396 2456 27402 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 36357 2459 36415 2465
rect 4387 2400 5580 2428
rect 7009 2431 7067 2437
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8294 2428 8300 2440
rect 7055 2400 8300 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 15010 2388 15016 2440
rect 15068 2388 15074 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22060 2400 22661 2428
rect 22060 2388 22066 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25464 2400 25697 2428
rect 25464 2388 25470 2400
rect 25685 2397 25697 2400
rect 25731 2428 25743 2431
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25731 2400 25973 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33468 2400 33701 2428
rect 33468 2388 33474 2400
rect 33689 2397 33701 2400
rect 33735 2428 33747 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33735 2400 33977 2428
rect 33735 2397 33747 2400
rect 33689 2391 33747 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36136 2400 37289 2428
rect 36136 2388 36142 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 4890 2360 4896 2372
rect 1872 2332 4896 2360
rect 4890 2320 4896 2332
rect 4948 2320 4954 2372
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 22836 25644 22888 25696
rect 27804 25644 27856 25696
rect 10140 25576 10192 25628
rect 33600 25576 33652 25628
rect 7012 25508 7064 25560
rect 32864 25508 32916 25560
rect 10876 25440 10928 25492
rect 35624 25440 35676 25492
rect 15844 25372 15896 25424
rect 34244 25372 34296 25424
rect 10048 25304 10100 25356
rect 31576 25304 31628 25356
rect 12072 25236 12124 25288
rect 33784 25236 33836 25288
rect 12624 25168 12676 25220
rect 34796 25168 34848 25220
rect 9864 25100 9916 25152
rect 31760 25100 31812 25152
rect 10784 25032 10836 25084
rect 34612 25032 34664 25084
rect 14924 24964 14976 25016
rect 31116 24964 31168 25016
rect 4068 24896 4120 24948
rect 7472 24896 7524 24948
rect 15384 24896 15436 24948
rect 33692 24896 33744 24948
rect 12808 24828 12860 24880
rect 32036 24828 32088 24880
rect 11704 24760 11756 24812
rect 22008 24760 22060 24812
rect 22560 24760 22612 24812
rect 30012 24760 30064 24812
rect 14280 24692 14332 24744
rect 26056 24692 26108 24744
rect 12348 24624 12400 24676
rect 25780 24624 25832 24676
rect 25964 24624 26016 24676
rect 30380 24692 30432 24744
rect 28264 24624 28316 24676
rect 31208 24624 31260 24676
rect 35900 24624 35952 24676
rect 36820 24624 36872 24676
rect 17132 24556 17184 24608
rect 18788 24556 18840 24608
rect 25136 24556 25188 24608
rect 29000 24556 29052 24608
rect 29092 24556 29144 24608
rect 40316 24556 40368 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 2044 24284 2096 24336
rect 3516 24216 3568 24268
rect 2320 24148 2372 24200
rect 4252 24148 4304 24200
rect 7104 24216 7156 24268
rect 9312 24284 9364 24336
rect 11704 24395 11756 24404
rect 11704 24361 11713 24395
rect 11713 24361 11747 24395
rect 11747 24361 11756 24395
rect 11704 24352 11756 24361
rect 14280 24395 14332 24404
rect 14280 24361 14289 24395
rect 14289 24361 14323 24395
rect 14323 24361 14332 24395
rect 14280 24352 14332 24361
rect 14464 24284 14516 24336
rect 6644 24148 6696 24200
rect 7196 24191 7248 24200
rect 7196 24157 7205 24191
rect 7205 24157 7239 24191
rect 7239 24157 7248 24191
rect 7196 24148 7248 24157
rect 3608 24012 3660 24064
rect 6000 24012 6052 24064
rect 6552 24055 6604 24064
rect 6552 24021 6561 24055
rect 6561 24021 6595 24055
rect 6595 24021 6604 24055
rect 6552 24012 6604 24021
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 10048 24148 10100 24200
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12624 24148 12676 24200
rect 18972 24352 19024 24404
rect 20168 24352 20220 24404
rect 41512 24352 41564 24404
rect 18144 24284 18196 24336
rect 18696 24216 18748 24268
rect 19064 24284 19116 24336
rect 13912 24148 13964 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 13820 24080 13872 24132
rect 19524 24148 19576 24200
rect 19892 24148 19944 24200
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21548 24216 21600 24268
rect 21180 24148 21232 24200
rect 22008 24191 22060 24200
rect 22008 24157 22017 24191
rect 22017 24157 22051 24191
rect 22051 24157 22060 24191
rect 22008 24148 22060 24157
rect 22100 24148 22152 24200
rect 25044 24216 25096 24268
rect 25136 24259 25188 24268
rect 25136 24225 25145 24259
rect 25145 24225 25179 24259
rect 25179 24225 25188 24259
rect 25136 24216 25188 24225
rect 25228 24216 25280 24268
rect 27620 24284 27672 24336
rect 28632 24216 28684 24268
rect 29276 24216 29328 24268
rect 33508 24327 33560 24336
rect 33508 24293 33517 24327
rect 33517 24293 33551 24327
rect 33551 24293 33560 24327
rect 33508 24284 33560 24293
rect 34060 24284 34112 24336
rect 34244 24259 34296 24268
rect 34244 24225 34253 24259
rect 34253 24225 34287 24259
rect 34287 24225 34296 24259
rect 34244 24216 34296 24225
rect 25320 24148 25372 24200
rect 17040 24080 17092 24132
rect 17132 24123 17184 24132
rect 17132 24089 17141 24123
rect 17141 24089 17175 24123
rect 17175 24089 17184 24123
rect 17132 24080 17184 24089
rect 18512 24080 18564 24132
rect 13728 24012 13780 24064
rect 16948 24012 17000 24064
rect 18788 24012 18840 24064
rect 25228 24080 25280 24132
rect 20444 24012 20496 24064
rect 24492 24012 24544 24064
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 24952 24055 25004 24064
rect 24952 24021 24961 24055
rect 24961 24021 24995 24055
rect 24995 24021 25004 24055
rect 24952 24012 25004 24021
rect 25964 24080 26016 24132
rect 26056 24080 26108 24132
rect 26700 24080 26752 24132
rect 29184 24191 29236 24200
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 30012 24191 30064 24200
rect 30012 24157 30021 24191
rect 30021 24157 30055 24191
rect 30055 24157 30064 24191
rect 30012 24148 30064 24157
rect 30564 24148 30616 24200
rect 31484 24191 31536 24200
rect 31484 24157 31493 24191
rect 31493 24157 31527 24191
rect 31527 24157 31536 24191
rect 31484 24148 31536 24157
rect 31852 24148 31904 24200
rect 32496 24191 32548 24200
rect 32496 24157 32505 24191
rect 32505 24157 32539 24191
rect 32539 24157 32548 24191
rect 32496 24148 32548 24157
rect 33324 24191 33376 24200
rect 33324 24157 33333 24191
rect 33333 24157 33367 24191
rect 33367 24157 33376 24191
rect 33324 24148 33376 24157
rect 34060 24191 34112 24200
rect 34060 24157 34069 24191
rect 34069 24157 34103 24191
rect 34103 24157 34112 24191
rect 34060 24148 34112 24157
rect 34520 24148 34572 24200
rect 39580 24216 39632 24268
rect 40316 24259 40368 24268
rect 40316 24225 40325 24259
rect 40325 24225 40359 24259
rect 40359 24225 40368 24259
rect 40316 24216 40368 24225
rect 35072 24148 35124 24200
rect 30932 24080 30984 24132
rect 25780 24055 25832 24064
rect 25780 24021 25789 24055
rect 25789 24021 25823 24055
rect 25823 24021 25832 24055
rect 25780 24012 25832 24021
rect 26148 24055 26200 24064
rect 26148 24021 26157 24055
rect 26157 24021 26191 24055
rect 26191 24021 26200 24055
rect 26148 24012 26200 24021
rect 27160 24055 27212 24064
rect 27160 24021 27169 24055
rect 27169 24021 27203 24055
rect 27203 24021 27212 24055
rect 27160 24012 27212 24021
rect 27252 24012 27304 24064
rect 28356 24055 28408 24064
rect 28356 24021 28365 24055
rect 28365 24021 28399 24055
rect 28399 24021 28408 24055
rect 28356 24012 28408 24021
rect 29552 24012 29604 24064
rect 31392 24012 31444 24064
rect 31852 24012 31904 24064
rect 34612 24012 34664 24064
rect 36820 24148 36872 24200
rect 37280 24148 37332 24200
rect 38476 24191 38528 24200
rect 38476 24157 38485 24191
rect 38485 24157 38519 24191
rect 38519 24157 38528 24191
rect 38476 24148 38528 24157
rect 39212 24191 39264 24200
rect 39212 24157 39221 24191
rect 39221 24157 39255 24191
rect 39255 24157 39264 24191
rect 39212 24148 39264 24157
rect 40592 24148 40644 24200
rect 44732 24395 44784 24404
rect 44732 24361 44741 24395
rect 44741 24361 44775 24395
rect 44775 24361 44784 24395
rect 44732 24352 44784 24361
rect 44732 24148 44784 24200
rect 45284 24148 45336 24200
rect 35900 24123 35952 24132
rect 35900 24089 35909 24123
rect 35909 24089 35943 24123
rect 35943 24089 35952 24123
rect 35900 24080 35952 24089
rect 40040 24080 40092 24132
rect 45560 24148 45612 24200
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 47952 24148 48004 24200
rect 36176 24012 36228 24064
rect 37464 24055 37516 24064
rect 37464 24021 37473 24055
rect 37473 24021 37507 24055
rect 37507 24021 37516 24055
rect 37464 24012 37516 24021
rect 39304 24055 39356 24064
rect 39304 24021 39313 24055
rect 39313 24021 39347 24055
rect 39347 24021 39356 24055
rect 39304 24012 39356 24021
rect 41328 24055 41380 24064
rect 41328 24021 41337 24055
rect 41337 24021 41371 24055
rect 41371 24021 41380 24055
rect 41328 24012 41380 24021
rect 43996 24012 44048 24064
rect 45468 24012 45520 24064
rect 46848 24055 46900 24064
rect 46848 24021 46857 24055
rect 46857 24021 46891 24055
rect 46891 24021 46900 24055
rect 46848 24012 46900 24021
rect 48688 24055 48740 24064
rect 48688 24021 48697 24055
rect 48697 24021 48731 24055
rect 48731 24021 48740 24055
rect 48688 24012 48740 24021
rect 49516 24055 49568 24064
rect 49516 24021 49525 24055
rect 49525 24021 49559 24055
rect 49559 24021 49568 24055
rect 49516 24012 49568 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 3516 23808 3568 23860
rect 4988 23808 5040 23860
rect 4160 23740 4212 23792
rect 2596 23672 2648 23724
rect 3792 23672 3844 23724
rect 7288 23740 7340 23792
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 4068 23536 4120 23588
rect 6920 23604 6972 23656
rect 5908 23536 5960 23588
rect 7564 23604 7616 23656
rect 12348 23851 12400 23860
rect 12348 23817 12357 23851
rect 12357 23817 12391 23851
rect 12391 23817 12400 23851
rect 12348 23808 12400 23817
rect 17960 23808 18012 23860
rect 21180 23808 21232 23860
rect 9956 23740 10008 23792
rect 12532 23740 12584 23792
rect 15752 23740 15804 23792
rect 18328 23740 18380 23792
rect 19064 23740 19116 23792
rect 20720 23740 20772 23792
rect 22744 23740 22796 23792
rect 24952 23808 25004 23860
rect 27160 23808 27212 23860
rect 27712 23808 27764 23860
rect 25596 23740 25648 23792
rect 28172 23740 28224 23792
rect 8760 23672 8812 23724
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 12256 23715 12308 23724
rect 12256 23681 12265 23715
rect 12265 23681 12299 23715
rect 12299 23681 12308 23715
rect 12256 23672 12308 23681
rect 12624 23672 12676 23724
rect 14280 23672 14332 23724
rect 18144 23672 18196 23724
rect 18696 23715 18748 23724
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 1768 23468 1820 23520
rect 2780 23468 2832 23520
rect 5264 23468 5316 23520
rect 6184 23468 6236 23520
rect 6736 23511 6788 23520
rect 6736 23477 6745 23511
rect 6745 23477 6779 23511
rect 6779 23477 6788 23511
rect 6736 23468 6788 23477
rect 6920 23468 6972 23520
rect 7748 23468 7800 23520
rect 11520 23511 11572 23520
rect 11520 23477 11529 23511
rect 11529 23477 11563 23511
rect 11563 23477 11572 23511
rect 11520 23468 11572 23477
rect 11888 23511 11940 23520
rect 11888 23477 11897 23511
rect 11897 23477 11931 23511
rect 11931 23477 11940 23511
rect 11888 23468 11940 23477
rect 16948 23604 17000 23656
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 19340 23604 19392 23656
rect 29552 23715 29604 23724
rect 29552 23681 29561 23715
rect 29561 23681 29595 23715
rect 29595 23681 29604 23715
rect 29552 23672 29604 23681
rect 30932 23851 30984 23860
rect 30932 23817 30941 23851
rect 30941 23817 30975 23851
rect 30975 23817 30984 23851
rect 30932 23808 30984 23817
rect 31116 23808 31168 23860
rect 32864 23808 32916 23860
rect 33600 23808 33652 23860
rect 34796 23851 34848 23860
rect 34796 23817 34805 23851
rect 34805 23817 34839 23851
rect 34839 23817 34848 23851
rect 34796 23808 34848 23817
rect 34980 23808 35032 23860
rect 37464 23808 37516 23860
rect 38476 23851 38528 23860
rect 38476 23817 38485 23851
rect 38485 23817 38519 23851
rect 38519 23817 38528 23851
rect 38476 23808 38528 23817
rect 39212 23808 39264 23860
rect 39580 23808 39632 23860
rect 43444 23808 43496 23860
rect 45560 23808 45612 23860
rect 47308 23808 47360 23860
rect 30104 23783 30156 23792
rect 30104 23749 30113 23783
rect 30113 23749 30147 23783
rect 30147 23749 30156 23783
rect 30104 23740 30156 23749
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 23296 23604 23348 23656
rect 24400 23536 24452 23588
rect 15108 23468 15160 23520
rect 18696 23468 18748 23520
rect 20076 23468 20128 23520
rect 20536 23468 20588 23520
rect 23848 23468 23900 23520
rect 24584 23468 24636 23520
rect 25136 23647 25188 23656
rect 25136 23613 25145 23647
rect 25145 23613 25179 23647
rect 25179 23613 25188 23647
rect 25136 23604 25188 23613
rect 27160 23647 27212 23656
rect 25688 23468 25740 23520
rect 27160 23613 27169 23647
rect 27169 23613 27203 23647
rect 27203 23613 27212 23647
rect 27160 23604 27212 23613
rect 27528 23604 27580 23656
rect 30932 23604 30984 23656
rect 31208 23672 31260 23724
rect 32588 23672 32640 23724
rect 35624 23783 35676 23792
rect 35624 23749 35633 23783
rect 35633 23749 35667 23783
rect 35667 23749 35676 23783
rect 35624 23740 35676 23749
rect 31852 23604 31904 23656
rect 26240 23468 26292 23520
rect 28448 23536 28500 23588
rect 28724 23468 28776 23520
rect 29184 23468 29236 23520
rect 32128 23579 32180 23588
rect 32128 23545 32137 23579
rect 32137 23545 32171 23579
rect 32171 23545 32180 23579
rect 32404 23604 32456 23656
rect 34888 23672 34940 23724
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 36360 23672 36412 23724
rect 37648 23672 37700 23724
rect 41144 23672 41196 23724
rect 44180 23672 44232 23724
rect 46664 23672 46716 23724
rect 48320 23715 48372 23724
rect 48320 23681 48329 23715
rect 48329 23681 48363 23715
rect 48363 23681 48372 23715
rect 48320 23672 48372 23681
rect 49516 23672 49568 23724
rect 34612 23604 34664 23656
rect 32128 23536 32180 23545
rect 34704 23536 34756 23588
rect 41604 23604 41656 23656
rect 45468 23604 45520 23656
rect 29552 23468 29604 23520
rect 30472 23468 30524 23520
rect 36084 23511 36136 23520
rect 36084 23477 36093 23511
rect 36093 23477 36127 23511
rect 36127 23477 36136 23511
rect 36084 23468 36136 23477
rect 36728 23511 36780 23520
rect 36728 23477 36737 23511
rect 36737 23477 36771 23511
rect 36771 23477 36780 23511
rect 36728 23468 36780 23477
rect 41420 23468 41472 23520
rect 44456 23511 44508 23520
rect 44456 23477 44465 23511
rect 44465 23477 44499 23511
rect 44499 23477 44508 23511
rect 44456 23468 44508 23477
rect 46940 23511 46992 23520
rect 46940 23477 46949 23511
rect 46949 23477 46983 23511
rect 46983 23477 46992 23511
rect 46940 23468 46992 23477
rect 48504 23511 48556 23520
rect 48504 23477 48513 23511
rect 48513 23477 48547 23511
rect 48547 23477 48556 23511
rect 48504 23468 48556 23477
rect 49240 23511 49292 23520
rect 49240 23477 49249 23511
rect 49249 23477 49283 23511
rect 49283 23477 49292 23511
rect 49240 23468 49292 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 1860 23264 1912 23316
rect 17868 23264 17920 23316
rect 19616 23264 19668 23316
rect 19708 23264 19760 23316
rect 22100 23264 22152 23316
rect 22192 23264 22244 23316
rect 24308 23264 24360 23316
rect 24400 23264 24452 23316
rect 5172 23196 5224 23248
rect 13728 23196 13780 23248
rect 16580 23196 16632 23248
rect 19064 23196 19116 23248
rect 2872 23128 2924 23180
rect 4344 23128 4396 23180
rect 4804 23171 4856 23180
rect 4804 23137 4813 23171
rect 4813 23137 4847 23171
rect 4847 23137 4856 23171
rect 4804 23128 4856 23137
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 12440 23128 12492 23180
rect 17408 23128 17460 23180
rect 1952 23060 2004 23112
rect 4160 23060 4212 23112
rect 4528 23060 4580 23112
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 3976 22992 4028 23044
rect 6276 23060 6328 23112
rect 8300 23060 8352 23112
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 16856 23060 16908 23112
rect 18512 23060 18564 23112
rect 8484 22992 8536 23044
rect 3700 22924 3752 22976
rect 4712 22924 4764 22976
rect 9036 22967 9088 22976
rect 9036 22933 9045 22967
rect 9045 22933 9079 22967
rect 9079 22933 9088 22967
rect 9036 22924 9088 22933
rect 9588 23035 9640 23044
rect 9588 23001 9597 23035
rect 9597 23001 9631 23035
rect 9631 23001 9640 23035
rect 9588 22992 9640 23001
rect 11152 22992 11204 23044
rect 11520 22992 11572 23044
rect 11888 22992 11940 23044
rect 13176 22992 13228 23044
rect 13820 23035 13872 23044
rect 13820 23001 13829 23035
rect 13829 23001 13863 23035
rect 13863 23001 13872 23035
rect 13820 22992 13872 23001
rect 14372 23035 14424 23044
rect 14372 23001 14381 23035
rect 14381 23001 14415 23035
rect 14415 23001 14424 23035
rect 14372 22992 14424 23001
rect 16948 22992 17000 23044
rect 13452 22924 13504 22976
rect 16672 22924 16724 22976
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 22284 23196 22336 23248
rect 24308 23128 24360 23180
rect 19800 23060 19852 23112
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 24124 23060 24176 23112
rect 28724 23264 28776 23316
rect 29000 23307 29052 23316
rect 29000 23273 29009 23307
rect 29009 23273 29043 23307
rect 29043 23273 29052 23307
rect 29000 23264 29052 23273
rect 31208 23264 31260 23316
rect 32036 23264 32088 23316
rect 32680 23264 32732 23316
rect 36268 23264 36320 23316
rect 36820 23307 36872 23316
rect 36820 23273 36829 23307
rect 36829 23273 36863 23307
rect 36863 23273 36872 23307
rect 36820 23264 36872 23273
rect 37280 23307 37332 23316
rect 37280 23273 37289 23307
rect 37289 23273 37323 23307
rect 37323 23273 37332 23307
rect 37280 23264 37332 23273
rect 27160 23128 27212 23180
rect 28540 23196 28592 23248
rect 27620 23128 27672 23180
rect 28172 23128 28224 23180
rect 29092 23128 29144 23180
rect 31484 23196 31536 23248
rect 35992 23239 36044 23248
rect 35992 23205 36001 23239
rect 36001 23205 36035 23239
rect 36035 23205 36044 23239
rect 35992 23196 36044 23205
rect 20352 23035 20404 23044
rect 20352 23001 20361 23035
rect 20361 23001 20395 23035
rect 20395 23001 20404 23035
rect 20352 22992 20404 23001
rect 20812 22992 20864 23044
rect 22836 22992 22888 23044
rect 20628 22924 20680 22976
rect 24768 22992 24820 23044
rect 25596 22992 25648 23044
rect 23296 22924 23348 22976
rect 23388 22924 23440 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 24952 22924 25004 22933
rect 26148 22967 26200 22976
rect 26148 22933 26157 22967
rect 26157 22933 26191 22967
rect 26191 22933 26200 22967
rect 26148 22924 26200 22933
rect 26516 22924 26568 22976
rect 28172 22992 28224 23044
rect 37832 23128 37884 23180
rect 33692 23060 33744 23112
rect 33784 23060 33836 23112
rect 34428 23060 34480 23112
rect 35716 23103 35768 23112
rect 35716 23069 35725 23103
rect 35725 23069 35759 23103
rect 35759 23069 35768 23103
rect 35716 23060 35768 23069
rect 35992 23060 36044 23112
rect 48596 23103 48648 23112
rect 48596 23069 48605 23103
rect 48605 23069 48639 23103
rect 48639 23069 48648 23103
rect 48596 23060 48648 23069
rect 49332 23060 49384 23112
rect 30012 22992 30064 23044
rect 30472 22992 30524 23044
rect 28356 22924 28408 22976
rect 29736 22924 29788 22976
rect 31484 22967 31536 22976
rect 31484 22933 31493 22967
rect 31493 22933 31527 22967
rect 31527 22933 31536 22967
rect 31484 22924 31536 22933
rect 31668 22924 31720 22976
rect 32128 22992 32180 23044
rect 33416 22992 33468 23044
rect 34520 22924 34572 22976
rect 35532 22967 35584 22976
rect 35532 22933 35541 22967
rect 35541 22933 35575 22967
rect 35575 22933 35584 22967
rect 35532 22924 35584 22933
rect 48412 22967 48464 22976
rect 48412 22933 48421 22967
rect 48421 22933 48455 22967
rect 48455 22933 48464 22967
rect 48412 22924 48464 22933
rect 48780 22924 48832 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 2228 22720 2280 22772
rect 4436 22720 4488 22772
rect 3700 22652 3752 22704
rect 1860 22584 1912 22636
rect 3608 22584 3660 22636
rect 4068 22652 4120 22704
rect 6920 22720 6972 22772
rect 9036 22720 9088 22772
rect 14464 22720 14516 22772
rect 19708 22720 19760 22772
rect 20352 22720 20404 22772
rect 22192 22720 22244 22772
rect 23664 22720 23716 22772
rect 5356 22652 5408 22704
rect 2872 22516 2924 22568
rect 3424 22516 3476 22568
rect 4068 22559 4120 22568
rect 4068 22525 4077 22559
rect 4077 22525 4111 22559
rect 4111 22525 4120 22559
rect 4068 22516 4120 22525
rect 2412 22448 2464 22500
rect 3976 22448 4028 22500
rect 6644 22584 6696 22636
rect 6736 22584 6788 22636
rect 7656 22584 7708 22636
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 11796 22695 11848 22704
rect 11796 22661 11805 22695
rect 11805 22661 11839 22695
rect 11839 22661 11848 22695
rect 11796 22652 11848 22661
rect 11888 22652 11940 22704
rect 13176 22652 13228 22704
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 17132 22695 17184 22704
rect 17132 22661 17141 22695
rect 17141 22661 17175 22695
rect 17175 22661 17184 22695
rect 17132 22652 17184 22661
rect 18512 22652 18564 22704
rect 10140 22584 10192 22636
rect 16764 22584 16816 22636
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19432 22584 19484 22636
rect 20076 22652 20128 22704
rect 20720 22652 20772 22704
rect 22284 22584 22336 22636
rect 23296 22652 23348 22704
rect 23388 22695 23440 22704
rect 23388 22661 23397 22695
rect 23397 22661 23431 22695
rect 23431 22661 23440 22695
rect 23388 22652 23440 22661
rect 23480 22652 23532 22704
rect 24676 22720 24728 22772
rect 25688 22720 25740 22772
rect 28448 22720 28500 22772
rect 25136 22652 25188 22704
rect 27344 22652 27396 22704
rect 24768 22584 24820 22636
rect 24952 22584 25004 22636
rect 27436 22584 27488 22636
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 7380 22559 7432 22568
rect 7380 22525 7389 22559
rect 7389 22525 7423 22559
rect 7423 22525 7432 22559
rect 7380 22516 7432 22525
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 13452 22516 13504 22568
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 3700 22380 3752 22432
rect 6368 22423 6420 22432
rect 6368 22389 6377 22423
rect 6377 22389 6411 22423
rect 6411 22389 6420 22423
rect 6368 22380 6420 22389
rect 6460 22380 6512 22432
rect 7104 22380 7156 22432
rect 16120 22448 16172 22500
rect 16212 22448 16264 22500
rect 20536 22516 20588 22568
rect 20628 22516 20680 22568
rect 23388 22516 23440 22568
rect 23940 22516 23992 22568
rect 27620 22559 27672 22568
rect 27620 22525 27629 22559
rect 27629 22525 27663 22559
rect 27663 22525 27672 22559
rect 27620 22516 27672 22525
rect 28540 22652 28592 22704
rect 31484 22720 31536 22772
rect 31760 22720 31812 22772
rect 33324 22720 33376 22772
rect 29092 22652 29144 22704
rect 36084 22652 36136 22704
rect 40040 22720 40092 22772
rect 48596 22720 48648 22772
rect 49332 22763 49384 22772
rect 49332 22729 49341 22763
rect 49341 22729 49375 22763
rect 49375 22729 49384 22763
rect 49332 22720 49384 22729
rect 31208 22584 31260 22636
rect 32864 22584 32916 22636
rect 32956 22584 33008 22636
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 37832 22627 37884 22636
rect 37832 22593 37841 22627
rect 37841 22593 37875 22627
rect 37875 22593 37884 22627
rect 37832 22584 37884 22593
rect 18788 22448 18840 22500
rect 14188 22423 14240 22432
rect 14188 22389 14197 22423
rect 14197 22389 14231 22423
rect 14231 22389 14240 22423
rect 14188 22380 14240 22389
rect 16764 22380 16816 22432
rect 18420 22380 18472 22432
rect 19156 22380 19208 22432
rect 21824 22380 21876 22432
rect 23480 22380 23532 22432
rect 25412 22448 25464 22500
rect 28724 22516 28776 22568
rect 30012 22448 30064 22500
rect 31668 22516 31720 22568
rect 33324 22516 33376 22568
rect 31300 22448 31352 22500
rect 35716 22448 35768 22500
rect 26516 22423 26568 22432
rect 26516 22389 26525 22423
rect 26525 22389 26559 22423
rect 26559 22389 26568 22423
rect 26516 22380 26568 22389
rect 28448 22380 28500 22432
rect 29092 22380 29144 22432
rect 30380 22380 30432 22432
rect 32864 22423 32916 22432
rect 32864 22389 32873 22423
rect 32873 22389 32907 22423
rect 32907 22389 32916 22423
rect 32864 22380 32916 22389
rect 33416 22380 33468 22432
rect 34520 22380 34572 22432
rect 34888 22423 34940 22432
rect 34888 22389 34897 22423
rect 34897 22389 34931 22423
rect 34931 22389 34940 22423
rect 34888 22380 34940 22389
rect 48412 22516 48464 22568
rect 49516 22423 49568 22432
rect 49516 22389 49525 22423
rect 49525 22389 49559 22423
rect 49559 22389 49568 22423
rect 49516 22380 49568 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 1952 22176 2004 22228
rect 3976 22108 4028 22160
rect 7104 22108 7156 22160
rect 9680 22108 9732 22160
rect 11980 22108 12032 22160
rect 12532 22108 12584 22160
rect 1308 22040 1360 22092
rect 3240 22040 3292 22092
rect 3976 21972 4028 22024
rect 8852 22040 8904 22092
rect 9220 22083 9272 22092
rect 9220 22049 9229 22083
rect 9229 22049 9263 22083
rect 9263 22049 9272 22083
rect 9220 22040 9272 22049
rect 10140 22040 10192 22092
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 15016 22176 15068 22228
rect 17132 22176 17184 22228
rect 18512 22108 18564 22160
rect 19064 22108 19116 22160
rect 19432 22040 19484 22092
rect 6552 21972 6604 22024
rect 7104 21972 7156 22024
rect 9496 21972 9548 22024
rect 10048 21972 10100 22024
rect 10784 21972 10836 22024
rect 12808 21972 12860 22024
rect 15016 21972 15068 22024
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 15384 21972 15436 21981
rect 18512 21972 18564 22024
rect 18880 21972 18932 22024
rect 25044 22176 25096 22228
rect 20260 22108 20312 22160
rect 24676 22108 24728 22160
rect 28816 22176 28868 22228
rect 34520 22176 34572 22228
rect 27068 22108 27120 22160
rect 26424 22040 26476 22092
rect 27344 22108 27396 22160
rect 31484 22108 31536 22160
rect 31668 22108 31720 22160
rect 40040 22176 40092 22228
rect 31576 22083 31628 22092
rect 31576 22049 31585 22083
rect 31585 22049 31619 22083
rect 31619 22049 31628 22083
rect 31576 22040 31628 22049
rect 32496 22040 32548 22092
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 25412 21972 25464 22024
rect 25596 21972 25648 22024
rect 27804 21972 27856 22024
rect 6828 21904 6880 21956
rect 11796 21904 11848 21956
rect 17500 21904 17552 21956
rect 3424 21836 3476 21888
rect 5816 21879 5868 21888
rect 5816 21845 5825 21879
rect 5825 21845 5859 21879
rect 5859 21845 5868 21879
rect 5816 21836 5868 21845
rect 6092 21879 6144 21888
rect 6092 21845 6101 21879
rect 6101 21845 6135 21879
rect 6135 21845 6144 21879
rect 6092 21836 6144 21845
rect 7748 21836 7800 21888
rect 8392 21836 8444 21888
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 9404 21836 9456 21888
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 11428 21836 11480 21888
rect 11520 21836 11572 21888
rect 19984 21947 20036 21956
rect 19984 21913 19993 21947
rect 19993 21913 20027 21947
rect 20027 21913 20036 21947
rect 19984 21904 20036 21913
rect 21364 21904 21416 21956
rect 25228 21904 25280 21956
rect 26516 21904 26568 21956
rect 29000 21904 29052 21956
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 20076 21836 20128 21888
rect 21732 21836 21784 21888
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 22376 21836 22428 21888
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 23664 21836 23716 21845
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 27344 21836 27396 21888
rect 28356 21836 28408 21888
rect 28540 21836 28592 21888
rect 28632 21879 28684 21888
rect 28632 21845 28641 21879
rect 28641 21845 28675 21879
rect 28675 21845 28684 21879
rect 28632 21836 28684 21845
rect 29184 21879 29236 21888
rect 29184 21845 29193 21879
rect 29193 21845 29227 21879
rect 29227 21845 29236 21879
rect 29184 21836 29236 21845
rect 30012 21836 30064 21888
rect 30472 21947 30524 21956
rect 30472 21913 30481 21947
rect 30481 21913 30515 21947
rect 30515 21913 30524 21947
rect 30472 21904 30524 21913
rect 31300 21904 31352 21956
rect 32128 21972 32180 22024
rect 32772 21972 32824 22024
rect 49516 21972 49568 22024
rect 31024 21836 31076 21888
rect 36176 21904 36228 21956
rect 32036 21836 32088 21888
rect 48320 21836 48372 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 5540 21632 5592 21684
rect 4344 21607 4396 21616
rect 4344 21573 4353 21607
rect 4353 21573 4387 21607
rect 4387 21573 4396 21607
rect 4344 21564 4396 21573
rect 5816 21564 5868 21616
rect 7564 21564 7616 21616
rect 7840 21564 7892 21616
rect 8944 21564 8996 21616
rect 2228 21496 2280 21548
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 1400 21428 1452 21480
rect 2136 21360 2188 21412
rect 6644 21428 6696 21480
rect 4896 21360 4948 21412
rect 5540 21292 5592 21344
rect 6368 21335 6420 21344
rect 6368 21301 6377 21335
rect 6377 21301 6411 21335
rect 6411 21301 6420 21335
rect 6368 21292 6420 21301
rect 7012 21292 7064 21344
rect 9496 21632 9548 21684
rect 9772 21632 9824 21684
rect 12164 21632 12216 21684
rect 9588 21564 9640 21616
rect 9772 21496 9824 21548
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 11980 21496 12032 21548
rect 12348 21564 12400 21616
rect 14188 21632 14240 21684
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 17684 21632 17736 21684
rect 17776 21632 17828 21684
rect 20260 21632 20312 21684
rect 23480 21632 23532 21684
rect 13820 21564 13872 21616
rect 15384 21564 15436 21616
rect 18512 21564 18564 21616
rect 9864 21428 9916 21480
rect 12256 21471 12308 21480
rect 10232 21360 10284 21412
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 12440 21496 12492 21548
rect 15108 21496 15160 21548
rect 16672 21496 16724 21548
rect 17040 21539 17092 21548
rect 17040 21505 17049 21539
rect 17049 21505 17083 21539
rect 17083 21505 17092 21539
rect 17040 21496 17092 21505
rect 13452 21428 13504 21480
rect 14464 21360 14516 21412
rect 15292 21360 15344 21412
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 16212 21471 16264 21480
rect 16212 21437 16221 21471
rect 16221 21437 16255 21471
rect 16255 21437 16264 21471
rect 16212 21428 16264 21437
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17684 21360 17736 21412
rect 8300 21292 8352 21344
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 9772 21292 9824 21301
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 15016 21292 15068 21344
rect 15660 21292 15712 21344
rect 18604 21292 18656 21344
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 19064 21428 19116 21480
rect 20720 21564 20772 21616
rect 24584 21632 24636 21684
rect 27068 21632 27120 21684
rect 27344 21632 27396 21684
rect 35532 21632 35584 21684
rect 36544 21632 36596 21684
rect 46940 21632 46992 21684
rect 23940 21564 23992 21616
rect 25136 21564 25188 21616
rect 20352 21428 20404 21480
rect 23296 21496 23348 21548
rect 24768 21496 24820 21548
rect 25228 21496 25280 21548
rect 29000 21564 29052 21616
rect 29184 21564 29236 21616
rect 36728 21564 36780 21616
rect 28080 21496 28132 21548
rect 28356 21496 28408 21548
rect 30932 21496 30984 21548
rect 31760 21539 31812 21548
rect 31760 21505 31769 21539
rect 31769 21505 31803 21539
rect 31803 21505 31812 21539
rect 31760 21496 31812 21505
rect 32404 21539 32456 21548
rect 32404 21505 32413 21539
rect 32413 21505 32447 21539
rect 32447 21505 32456 21539
rect 32404 21496 32456 21505
rect 47860 21496 47912 21548
rect 24676 21428 24728 21480
rect 20812 21360 20864 21412
rect 27896 21471 27948 21480
rect 27896 21437 27905 21471
rect 27905 21437 27939 21471
rect 27939 21437 27948 21471
rect 27896 21428 27948 21437
rect 29092 21428 29144 21480
rect 19432 21292 19484 21344
rect 19708 21292 19760 21344
rect 20720 21335 20772 21344
rect 20720 21301 20729 21335
rect 20729 21301 20763 21335
rect 20763 21301 20772 21335
rect 20720 21292 20772 21301
rect 21824 21292 21876 21344
rect 23480 21292 23532 21344
rect 24216 21292 24268 21344
rect 24308 21292 24360 21344
rect 28908 21292 28960 21344
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 30288 21360 30340 21412
rect 32128 21360 32180 21412
rect 32680 21360 32732 21412
rect 48504 21360 48556 21412
rect 30656 21335 30708 21344
rect 30656 21301 30665 21335
rect 30665 21301 30699 21335
rect 30699 21301 30708 21335
rect 30656 21292 30708 21301
rect 30932 21292 30984 21344
rect 32496 21335 32548 21344
rect 32496 21301 32505 21335
rect 32505 21301 32539 21335
rect 32539 21301 32548 21335
rect 32496 21292 32548 21301
rect 47860 21292 47912 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 3424 21088 3476 21140
rect 7380 21088 7432 21140
rect 8576 21088 8628 21140
rect 8668 21088 8720 21140
rect 11520 21088 11572 21140
rect 3976 20995 4028 21004
rect 3976 20961 3985 20995
rect 3985 20961 4019 20995
rect 4019 20961 4028 20995
rect 3976 20952 4028 20961
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 7380 20952 7432 21004
rect 10600 21020 10652 21072
rect 11796 21020 11848 21072
rect 1860 20884 1912 20936
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 7012 20884 7064 20936
rect 8484 20995 8536 21004
rect 8484 20961 8493 20995
rect 8493 20961 8527 20995
rect 8527 20961 8536 20995
rect 8484 20952 8536 20961
rect 16028 21088 16080 21140
rect 16212 21088 16264 21140
rect 24124 21088 24176 21140
rect 12256 21020 12308 21072
rect 14096 21020 14148 21072
rect 2872 20816 2924 20868
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 12532 20952 12584 20961
rect 13820 20952 13872 21004
rect 14188 20995 14240 21004
rect 14188 20961 14197 20995
rect 14197 20961 14231 20995
rect 14231 20961 14240 20995
rect 14188 20952 14240 20961
rect 14464 20952 14516 21004
rect 15108 20995 15160 21004
rect 15108 20961 15117 20995
rect 15117 20961 15151 20995
rect 15151 20961 15160 20995
rect 15108 20952 15160 20961
rect 16764 21020 16816 21072
rect 11152 20884 11204 20936
rect 12072 20927 12124 20936
rect 12072 20893 12081 20927
rect 12081 20893 12115 20927
rect 12115 20893 12124 20927
rect 12072 20884 12124 20893
rect 16212 20927 16264 20936
rect 16212 20893 16221 20927
rect 16221 20893 16255 20927
rect 16255 20893 16264 20927
rect 16212 20884 16264 20893
rect 6368 20748 6420 20800
rect 8392 20816 8444 20868
rect 11336 20859 11388 20868
rect 11336 20825 11345 20859
rect 11345 20825 11379 20859
rect 11379 20825 11388 20859
rect 11336 20816 11388 20825
rect 7196 20791 7248 20800
rect 7196 20757 7205 20791
rect 7205 20757 7239 20791
rect 7239 20757 7248 20791
rect 7196 20748 7248 20757
rect 7380 20748 7432 20800
rect 8116 20748 8168 20800
rect 10600 20748 10652 20800
rect 11428 20791 11480 20800
rect 11428 20757 11437 20791
rect 11437 20757 11471 20791
rect 11471 20757 11480 20791
rect 11428 20748 11480 20757
rect 16488 20816 16540 20868
rect 17960 20952 18012 21004
rect 18788 20995 18840 21004
rect 18788 20961 18797 20995
rect 18797 20961 18831 20995
rect 18831 20961 18840 20995
rect 18788 20952 18840 20961
rect 21824 21063 21876 21072
rect 21824 21029 21833 21063
rect 21833 21029 21867 21063
rect 21867 21029 21876 21063
rect 21824 21020 21876 21029
rect 19708 20995 19760 21004
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 20260 20952 20312 21004
rect 24400 21020 24452 21072
rect 22744 20995 22796 21004
rect 22744 20961 22753 20995
rect 22753 20961 22787 20995
rect 22787 20961 22796 20995
rect 22744 20952 22796 20961
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 30656 21088 30708 21140
rect 32588 21088 32640 21140
rect 25964 21020 26016 21072
rect 27620 21020 27672 21072
rect 25596 20952 25648 21004
rect 26056 20995 26108 21004
rect 26056 20961 26065 20995
rect 26065 20961 26099 20995
rect 26099 20961 26108 20995
rect 26056 20952 26108 20961
rect 28356 20952 28408 21004
rect 28724 21020 28776 21072
rect 36544 21020 36596 21072
rect 30012 20995 30064 21004
rect 30012 20961 30021 20995
rect 30021 20961 30055 20995
rect 30055 20961 30064 20995
rect 30012 20952 30064 20961
rect 17408 20927 17460 20936
rect 17408 20893 17417 20927
rect 17417 20893 17451 20927
rect 17451 20893 17460 20927
rect 17408 20884 17460 20893
rect 18880 20884 18932 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 27620 20884 27672 20936
rect 15660 20748 15712 20800
rect 15752 20791 15804 20800
rect 15752 20757 15761 20791
rect 15761 20757 15795 20791
rect 15795 20757 15804 20791
rect 15752 20748 15804 20757
rect 16672 20748 16724 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17776 20748 17828 20800
rect 18328 20748 18380 20800
rect 20720 20816 20772 20868
rect 23388 20816 23440 20868
rect 23664 20859 23716 20868
rect 23664 20825 23673 20859
rect 23673 20825 23707 20859
rect 23707 20825 23716 20859
rect 23664 20816 23716 20825
rect 26240 20816 26292 20868
rect 20444 20748 20496 20800
rect 20536 20748 20588 20800
rect 22192 20748 22244 20800
rect 22560 20791 22612 20800
rect 22560 20757 22569 20791
rect 22569 20757 22603 20791
rect 22603 20757 22612 20791
rect 22560 20748 22612 20757
rect 22652 20748 22704 20800
rect 23480 20748 23532 20800
rect 24032 20748 24084 20800
rect 24768 20748 24820 20800
rect 25872 20748 25924 20800
rect 26608 20816 26660 20868
rect 28448 20884 28500 20936
rect 29000 20884 29052 20936
rect 27620 20748 27672 20800
rect 27988 20748 28040 20800
rect 28080 20748 28132 20800
rect 28816 20748 28868 20800
rect 30932 20816 30984 20868
rect 31116 20859 31168 20868
rect 31116 20825 31125 20859
rect 31125 20825 31159 20859
rect 31159 20825 31168 20859
rect 31116 20816 31168 20825
rect 31760 20816 31812 20868
rect 30380 20748 30432 20800
rect 31944 20791 31996 20800
rect 31944 20757 31953 20791
rect 31953 20757 31987 20791
rect 31987 20757 31996 20791
rect 31944 20748 31996 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 4344 20544 4396 20596
rect 11428 20544 11480 20596
rect 3884 20476 3936 20528
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 4068 20408 4120 20460
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 6092 20408 6144 20460
rect 6828 20340 6880 20392
rect 9956 20476 10008 20528
rect 11152 20476 11204 20528
rect 12532 20476 12584 20528
rect 13544 20476 13596 20528
rect 7380 20408 7432 20460
rect 8944 20408 8996 20460
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 12808 20408 12860 20460
rect 9404 20383 9456 20392
rect 9404 20349 9413 20383
rect 9413 20349 9447 20383
rect 9447 20349 9456 20383
rect 9404 20340 9456 20349
rect 9680 20383 9732 20392
rect 9680 20349 9689 20383
rect 9689 20349 9723 20383
rect 9723 20349 9732 20383
rect 9680 20340 9732 20349
rect 6092 20272 6144 20324
rect 7380 20272 7432 20324
rect 11152 20383 11204 20392
rect 11152 20349 11161 20383
rect 11161 20349 11195 20383
rect 11195 20349 11204 20383
rect 11152 20340 11204 20349
rect 12256 20340 12308 20392
rect 12532 20340 12584 20392
rect 13636 20408 13688 20460
rect 14464 20476 14516 20528
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 16948 20544 17000 20596
rect 18880 20587 18932 20596
rect 18880 20553 18889 20587
rect 18889 20553 18923 20587
rect 18923 20553 18932 20587
rect 18880 20544 18932 20553
rect 19064 20544 19116 20596
rect 19432 20544 19484 20596
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 13452 20272 13504 20324
rect 7104 20204 7156 20256
rect 9036 20204 9088 20256
rect 10140 20204 10192 20256
rect 10876 20204 10928 20256
rect 11888 20247 11940 20256
rect 11888 20213 11897 20247
rect 11897 20213 11931 20247
rect 11931 20213 11940 20247
rect 11888 20204 11940 20213
rect 12716 20204 12768 20256
rect 13636 20247 13688 20256
rect 13636 20213 13645 20247
rect 13645 20213 13679 20247
rect 13679 20213 13688 20247
rect 13636 20204 13688 20213
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 14648 20340 14700 20392
rect 17500 20408 17552 20460
rect 17132 20272 17184 20324
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 16764 20204 16816 20256
rect 17960 20340 18012 20392
rect 18880 20340 18932 20392
rect 19432 20408 19484 20460
rect 19616 20408 19668 20460
rect 20720 20476 20772 20528
rect 22008 20519 22060 20528
rect 22008 20485 22017 20519
rect 22017 20485 22051 20519
rect 22051 20485 22060 20519
rect 22008 20476 22060 20485
rect 23388 20587 23440 20596
rect 23388 20553 23397 20587
rect 23397 20553 23431 20587
rect 23431 20553 23440 20587
rect 23388 20544 23440 20553
rect 23664 20544 23716 20596
rect 24768 20544 24820 20596
rect 27252 20544 27304 20596
rect 25872 20476 25924 20528
rect 28540 20544 28592 20596
rect 34980 20544 35032 20596
rect 27804 20476 27856 20528
rect 28908 20476 28960 20528
rect 29092 20476 29144 20528
rect 23296 20408 23348 20460
rect 19616 20272 19668 20324
rect 17960 20204 18012 20256
rect 18696 20204 18748 20256
rect 18880 20204 18932 20256
rect 19248 20204 19300 20256
rect 20628 20340 20680 20392
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 24676 20340 24728 20392
rect 25136 20340 25188 20392
rect 26516 20408 26568 20460
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 25964 20340 26016 20392
rect 26332 20272 26384 20324
rect 22560 20204 22612 20256
rect 27436 20272 27488 20324
rect 30012 20340 30064 20392
rect 30196 20204 30248 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 4344 20000 4396 20052
rect 5448 20000 5500 20052
rect 6368 19864 6420 19916
rect 8300 20000 8352 20052
rect 9404 20000 9456 20052
rect 10876 20043 10928 20052
rect 10876 20009 10885 20043
rect 10885 20009 10919 20043
rect 10919 20009 10928 20043
rect 10876 20000 10928 20009
rect 11060 20000 11112 20052
rect 11796 20000 11848 20052
rect 13360 20000 13412 20052
rect 14004 20000 14056 20052
rect 15016 20000 15068 20052
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 19892 20000 19944 20052
rect 21180 20000 21232 20052
rect 23388 20000 23440 20052
rect 9036 19864 9088 19916
rect 12440 19932 12492 19984
rect 12808 19932 12860 19984
rect 14372 19932 14424 19984
rect 17776 19932 17828 19984
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 15476 19864 15528 19916
rect 18972 19864 19024 19916
rect 19248 19864 19300 19916
rect 10508 19796 10560 19848
rect 11060 19796 11112 19848
rect 12164 19839 12216 19848
rect 12164 19805 12173 19839
rect 12173 19805 12207 19839
rect 12207 19805 12216 19839
rect 12164 19796 12216 19805
rect 14464 19796 14516 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 18328 19796 18380 19848
rect 19064 19796 19116 19848
rect 2872 19728 2924 19780
rect 6184 19728 6236 19780
rect 7472 19728 7524 19780
rect 3700 19660 3752 19712
rect 4252 19660 4304 19712
rect 7840 19660 7892 19712
rect 8300 19660 8352 19712
rect 10968 19728 11020 19780
rect 12624 19728 12676 19780
rect 12808 19728 12860 19780
rect 11152 19660 11204 19712
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 12716 19660 12768 19712
rect 13636 19660 13688 19712
rect 13912 19703 13964 19712
rect 13912 19669 13921 19703
rect 13921 19669 13955 19703
rect 13955 19669 13964 19703
rect 13912 19660 13964 19669
rect 14188 19703 14240 19712
rect 14188 19669 14197 19703
rect 14197 19669 14231 19703
rect 14231 19669 14240 19703
rect 14188 19660 14240 19669
rect 14372 19660 14424 19712
rect 14832 19660 14884 19712
rect 15292 19728 15344 19780
rect 18972 19728 19024 19780
rect 20260 19932 20312 19984
rect 22928 19932 22980 19984
rect 19616 19864 19668 19916
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 23848 19907 23900 19916
rect 19708 19796 19760 19848
rect 19984 19728 20036 19780
rect 16396 19660 16448 19712
rect 16948 19660 17000 19712
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 18328 19660 18380 19712
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 19892 19660 19944 19712
rect 20720 19660 20772 19712
rect 21456 19660 21508 19712
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 27620 19975 27672 19984
rect 27620 19941 27629 19975
rect 27629 19941 27663 19975
rect 27663 19941 27672 19975
rect 27620 19932 27672 19941
rect 29736 19975 29788 19984
rect 29736 19941 29745 19975
rect 29745 19941 29779 19975
rect 29779 19941 29788 19975
rect 29736 19932 29788 19941
rect 30472 19975 30524 19984
rect 30472 19941 30481 19975
rect 30481 19941 30515 19975
rect 30515 19941 30524 19975
rect 30472 19932 30524 19941
rect 26148 19864 26200 19916
rect 27712 19864 27764 19916
rect 28632 19907 28684 19916
rect 28632 19873 28641 19907
rect 28641 19873 28675 19907
rect 28675 19873 28684 19907
rect 28632 19864 28684 19873
rect 48320 20000 48372 20052
rect 25504 19796 25556 19848
rect 25780 19796 25832 19848
rect 27528 19796 27580 19848
rect 31300 19907 31352 19916
rect 31300 19873 31309 19907
rect 31309 19873 31343 19907
rect 31343 19873 31352 19907
rect 31300 19864 31352 19873
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 24032 19728 24084 19780
rect 25228 19728 25280 19780
rect 25688 19728 25740 19780
rect 26608 19728 26660 19780
rect 28356 19728 28408 19780
rect 30472 19796 30524 19848
rect 34612 19796 34664 19848
rect 22284 19660 22336 19712
rect 23296 19703 23348 19712
rect 23296 19669 23305 19703
rect 23305 19669 23339 19703
rect 23339 19669 23348 19703
rect 23296 19660 23348 19669
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 27712 19660 27764 19712
rect 29092 19660 29144 19712
rect 30288 19703 30340 19712
rect 30288 19669 30297 19703
rect 30297 19669 30331 19703
rect 30331 19669 30340 19703
rect 30288 19660 30340 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 4896 19456 4948 19508
rect 3516 19388 3568 19440
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3700 19320 3752 19372
rect 4528 19320 4580 19372
rect 4896 19320 4948 19372
rect 6460 19456 6512 19508
rect 10324 19456 10376 19508
rect 10416 19499 10468 19508
rect 10416 19465 10425 19499
rect 10425 19465 10459 19499
rect 10459 19465 10468 19499
rect 10416 19456 10468 19465
rect 10968 19456 11020 19508
rect 14556 19456 14608 19508
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 6920 19388 6972 19440
rect 7564 19388 7616 19440
rect 9956 19388 10008 19440
rect 10692 19388 10744 19440
rect 6460 19320 6512 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 8668 19320 8720 19372
rect 11980 19388 12032 19440
rect 14188 19388 14240 19440
rect 7196 19252 7248 19304
rect 9680 19252 9732 19304
rect 11060 19252 11112 19304
rect 4528 19184 4580 19236
rect 13452 19295 13504 19304
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 13912 19252 13964 19304
rect 14372 19388 14424 19440
rect 14464 19388 14516 19440
rect 18512 19456 18564 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 19248 19456 19300 19508
rect 23296 19456 23348 19508
rect 23572 19456 23624 19508
rect 26240 19456 26292 19508
rect 26608 19456 26660 19508
rect 30380 19456 30432 19508
rect 15844 19320 15896 19372
rect 16028 19320 16080 19372
rect 14464 19252 14516 19304
rect 14832 19252 14884 19304
rect 15016 19252 15068 19304
rect 5448 19116 5500 19168
rect 6552 19116 6604 19168
rect 13268 19184 13320 19236
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 14372 19227 14424 19236
rect 14372 19193 14381 19227
rect 14381 19193 14415 19227
rect 14415 19193 14424 19227
rect 14372 19184 14424 19193
rect 16212 19252 16264 19304
rect 17776 19320 17828 19372
rect 17684 19252 17736 19304
rect 20076 19388 20128 19440
rect 20720 19388 20772 19440
rect 22652 19388 22704 19440
rect 23848 19388 23900 19440
rect 26332 19388 26384 19440
rect 29092 19388 29144 19440
rect 32312 19388 32364 19440
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18972 19320 19024 19372
rect 19064 19320 19116 19372
rect 22744 19320 22796 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 16488 19184 16540 19236
rect 16672 19184 16724 19236
rect 17500 19184 17552 19236
rect 15108 19116 15160 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 17684 19159 17736 19168
rect 17684 19125 17693 19159
rect 17693 19125 17727 19159
rect 17727 19125 17736 19159
rect 17684 19116 17736 19125
rect 18144 19252 18196 19304
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20628 19252 20680 19304
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 24860 19252 24912 19304
rect 18052 19184 18104 19236
rect 22008 19227 22060 19236
rect 22008 19193 22017 19227
rect 22017 19193 22051 19227
rect 22051 19193 22060 19227
rect 22008 19184 22060 19193
rect 22100 19184 22152 19236
rect 26516 19320 26568 19372
rect 27160 19320 27212 19372
rect 27712 19320 27764 19372
rect 30656 19363 30708 19372
rect 30656 19329 30665 19363
rect 30665 19329 30699 19363
rect 30699 19329 30708 19363
rect 30656 19320 30708 19329
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 27896 19252 27948 19304
rect 18788 19116 18840 19168
rect 20996 19116 21048 19168
rect 21088 19116 21140 19168
rect 22928 19116 22980 19168
rect 25320 19184 25372 19236
rect 27804 19116 27856 19168
rect 28356 19116 28408 19168
rect 28632 19116 28684 19168
rect 30012 19159 30064 19168
rect 30012 19125 30021 19159
rect 30021 19125 30055 19159
rect 30055 19125 30064 19159
rect 30012 19116 30064 19125
rect 30288 19116 30340 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 3976 18912 4028 18964
rect 5356 18912 5408 18964
rect 7564 18912 7616 18964
rect 7840 18912 7892 18964
rect 8116 18844 8168 18896
rect 11612 18955 11664 18964
rect 11612 18921 11621 18955
rect 11621 18921 11655 18955
rect 11655 18921 11664 18955
rect 11612 18912 11664 18921
rect 10508 18887 10560 18896
rect 10508 18853 10517 18887
rect 10517 18853 10551 18887
rect 10551 18853 10560 18887
rect 10508 18844 10560 18853
rect 1400 18776 1452 18828
rect 8484 18776 8536 18828
rect 8760 18776 8812 18828
rect 9036 18776 9088 18828
rect 10048 18819 10100 18828
rect 10048 18785 10057 18819
rect 10057 18785 10091 18819
rect 10091 18785 10100 18819
rect 10048 18776 10100 18785
rect 14832 18912 14884 18964
rect 12348 18844 12400 18896
rect 14372 18844 14424 18896
rect 12256 18819 12308 18828
rect 12256 18785 12265 18819
rect 12265 18785 12299 18819
rect 12299 18785 12308 18819
rect 12256 18776 12308 18785
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 13728 18776 13780 18828
rect 15016 18819 15068 18828
rect 15016 18785 15025 18819
rect 15025 18785 15059 18819
rect 15059 18785 15068 18819
rect 15016 18776 15068 18785
rect 4528 18708 4580 18760
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 10140 18708 10192 18760
rect 11796 18708 11848 18760
rect 14924 18708 14976 18760
rect 3884 18572 3936 18624
rect 3976 18615 4028 18624
rect 3976 18581 3985 18615
rect 3985 18581 4019 18615
rect 4019 18581 4028 18615
rect 3976 18572 4028 18581
rect 4804 18640 4856 18692
rect 6184 18572 6236 18624
rect 6368 18615 6420 18624
rect 6368 18581 6377 18615
rect 6377 18581 6411 18615
rect 6411 18581 6420 18615
rect 8760 18640 8812 18692
rect 6368 18572 6420 18581
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 9956 18640 10008 18692
rect 10232 18640 10284 18692
rect 8576 18572 8628 18581
rect 10416 18572 10468 18624
rect 11336 18572 11388 18624
rect 12992 18572 13044 18624
rect 13268 18572 13320 18624
rect 13728 18572 13780 18624
rect 22008 18912 22060 18964
rect 22652 18912 22704 18964
rect 23388 18955 23440 18964
rect 23388 18921 23397 18955
rect 23397 18921 23431 18955
rect 23431 18921 23440 18955
rect 23388 18912 23440 18921
rect 23848 18912 23900 18964
rect 24032 18955 24084 18964
rect 24032 18921 24041 18955
rect 24041 18921 24075 18955
rect 24075 18921 24084 18955
rect 25136 18955 25188 18964
rect 24032 18912 24084 18921
rect 25136 18921 25145 18955
rect 25145 18921 25179 18955
rect 25179 18921 25188 18955
rect 25136 18912 25188 18921
rect 25688 18912 25740 18964
rect 29092 18912 29144 18964
rect 30288 18912 30340 18964
rect 16488 18844 16540 18896
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 18328 18844 18380 18896
rect 20168 18844 20220 18896
rect 21088 18844 21140 18896
rect 26700 18844 26752 18896
rect 32680 18844 32732 18896
rect 19708 18776 19760 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 22008 18776 22060 18828
rect 16856 18708 16908 18760
rect 17132 18708 17184 18760
rect 18052 18708 18104 18760
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 18788 18708 18840 18760
rect 15476 18683 15528 18692
rect 15476 18649 15492 18683
rect 15492 18649 15526 18683
rect 15526 18649 15528 18683
rect 15476 18640 15528 18649
rect 15016 18572 15068 18624
rect 16212 18640 16264 18692
rect 16396 18572 16448 18624
rect 20076 18640 20128 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 18696 18572 18748 18624
rect 20260 18572 20312 18624
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 23664 18776 23716 18828
rect 25780 18776 25832 18828
rect 26148 18776 26200 18828
rect 28724 18776 28776 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 26792 18708 26844 18760
rect 27160 18708 27212 18760
rect 27620 18751 27672 18760
rect 27620 18717 27629 18751
rect 27629 18717 27663 18751
rect 27663 18717 27672 18751
rect 27620 18708 27672 18717
rect 28908 18708 28960 18760
rect 29828 18708 29880 18760
rect 22100 18572 22152 18624
rect 22468 18572 22520 18624
rect 24032 18572 24084 18624
rect 24216 18615 24268 18624
rect 24216 18581 24225 18615
rect 24225 18581 24259 18615
rect 24259 18581 24268 18615
rect 24216 18572 24268 18581
rect 25964 18640 26016 18692
rect 30748 18640 30800 18692
rect 29736 18615 29788 18624
rect 29736 18581 29745 18615
rect 29745 18581 29779 18615
rect 29779 18581 29788 18615
rect 29736 18572 29788 18581
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 3976 18368 4028 18420
rect 14648 18368 14700 18420
rect 15108 18368 15160 18420
rect 16488 18411 16540 18420
rect 16488 18377 16497 18411
rect 16497 18377 16531 18411
rect 16531 18377 16540 18411
rect 16488 18368 16540 18377
rect 20996 18368 21048 18420
rect 26792 18411 26844 18420
rect 26792 18377 26801 18411
rect 26801 18377 26835 18411
rect 26835 18377 26844 18411
rect 26792 18368 26844 18377
rect 30104 18368 30156 18420
rect 30840 18368 30892 18420
rect 33324 18368 33376 18420
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 4436 18343 4488 18352
rect 4436 18309 4445 18343
rect 4445 18309 4479 18343
rect 4479 18309 4488 18343
rect 4436 18300 4488 18309
rect 7196 18300 7248 18352
rect 9772 18343 9824 18352
rect 9772 18309 9781 18343
rect 9781 18309 9815 18343
rect 9815 18309 9824 18343
rect 9772 18300 9824 18309
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 6276 18232 6328 18284
rect 6920 18232 6972 18284
rect 5356 18164 5408 18216
rect 6000 18164 6052 18216
rect 7380 18096 7432 18148
rect 10508 18232 10560 18284
rect 8576 18164 8628 18216
rect 9588 18164 9640 18216
rect 14004 18300 14056 18352
rect 14556 18300 14608 18352
rect 14832 18300 14884 18352
rect 11888 18232 11940 18284
rect 12624 18232 12676 18284
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13544 18232 13596 18284
rect 14924 18232 14976 18284
rect 15016 18232 15068 18284
rect 15568 18232 15620 18284
rect 12256 18164 12308 18216
rect 9128 18096 9180 18148
rect 11612 18096 11664 18148
rect 11796 18096 11848 18148
rect 6828 18028 6880 18080
rect 6920 18028 6972 18080
rect 10232 18028 10284 18080
rect 12164 18028 12216 18080
rect 12716 18096 12768 18148
rect 13268 18139 13320 18148
rect 13268 18105 13277 18139
rect 13277 18105 13311 18139
rect 13311 18105 13320 18139
rect 13268 18096 13320 18105
rect 16948 18164 17000 18216
rect 17040 18164 17092 18216
rect 20168 18300 20220 18352
rect 22836 18343 22888 18352
rect 17592 18232 17644 18284
rect 19432 18232 19484 18284
rect 20260 18232 20312 18284
rect 20536 18232 20588 18284
rect 19616 18164 19668 18216
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20996 18096 21048 18148
rect 22836 18309 22845 18343
rect 22845 18309 22879 18343
rect 22879 18309 22888 18343
rect 22836 18300 22888 18309
rect 24032 18300 24084 18352
rect 25320 18343 25372 18352
rect 25320 18309 25329 18343
rect 25329 18309 25363 18343
rect 25363 18309 25372 18343
rect 25320 18300 25372 18309
rect 26056 18343 26108 18352
rect 26056 18309 26065 18343
rect 26065 18309 26099 18343
rect 26099 18309 26108 18343
rect 26056 18300 26108 18309
rect 28632 18300 28684 18352
rect 29092 18300 29144 18352
rect 21180 18275 21232 18284
rect 21180 18241 21189 18275
rect 21189 18241 21223 18275
rect 21223 18241 21232 18275
rect 21180 18232 21232 18241
rect 27804 18232 27856 18284
rect 30656 18275 30708 18284
rect 30656 18241 30665 18275
rect 30665 18241 30699 18275
rect 30699 18241 30708 18275
rect 30656 18232 30708 18241
rect 12808 18028 12860 18080
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 17684 18028 17736 18080
rect 20628 18028 20680 18080
rect 21916 18164 21968 18216
rect 21824 18028 21876 18080
rect 22468 18028 22520 18080
rect 26240 18164 26292 18216
rect 27068 18164 27120 18216
rect 30748 18207 30800 18216
rect 30748 18173 30757 18207
rect 30757 18173 30791 18207
rect 30791 18173 30800 18207
rect 30748 18164 30800 18173
rect 30840 18207 30892 18216
rect 30840 18173 30849 18207
rect 30849 18173 30883 18207
rect 30883 18173 30892 18207
rect 30840 18164 30892 18173
rect 41604 18232 41656 18284
rect 30380 18096 30432 18148
rect 24676 18028 24728 18080
rect 27344 18028 27396 18080
rect 29828 18071 29880 18080
rect 29828 18037 29837 18071
rect 29837 18037 29871 18071
rect 29871 18037 29880 18071
rect 29828 18028 29880 18037
rect 30748 18028 30800 18080
rect 41420 18028 41472 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 3608 17867 3660 17876
rect 3608 17833 3617 17867
rect 3617 17833 3651 17867
rect 3651 17833 3660 17867
rect 3608 17824 3660 17833
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 4804 17824 4856 17876
rect 7656 17824 7708 17876
rect 10324 17824 10376 17876
rect 11612 17867 11664 17876
rect 11612 17833 11621 17867
rect 11621 17833 11655 17867
rect 11655 17833 11664 17867
rect 11612 17824 11664 17833
rect 13360 17824 13412 17876
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 1860 17756 1912 17808
rect 7932 17756 7984 17808
rect 7840 17688 7892 17740
rect 4160 17620 4212 17672
rect 4620 17620 4672 17672
rect 7104 17620 7156 17672
rect 9404 17688 9456 17740
rect 9956 17688 10008 17740
rect 13268 17756 13320 17808
rect 14372 17756 14424 17808
rect 16120 17688 16172 17740
rect 17132 17824 17184 17876
rect 17316 17824 17368 17876
rect 21824 17867 21876 17876
rect 21824 17833 21833 17867
rect 21833 17833 21867 17867
rect 21867 17833 21876 17867
rect 21824 17824 21876 17833
rect 21916 17824 21968 17876
rect 27528 17824 27580 17876
rect 28632 17824 28684 17876
rect 28816 17824 28868 17876
rect 17592 17756 17644 17808
rect 21088 17756 21140 17808
rect 22008 17756 22060 17808
rect 26240 17756 26292 17808
rect 28448 17756 28500 17808
rect 16948 17688 17000 17740
rect 17224 17688 17276 17740
rect 20352 17688 20404 17740
rect 24584 17688 24636 17740
rect 24676 17688 24728 17740
rect 27804 17688 27856 17740
rect 1216 17552 1268 17604
rect 4344 17552 4396 17604
rect 6184 17552 6236 17604
rect 7472 17552 7524 17604
rect 7564 17552 7616 17604
rect 10232 17620 10284 17672
rect 10876 17620 10928 17672
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 9128 17595 9180 17604
rect 9128 17561 9137 17595
rect 9137 17561 9171 17595
rect 9171 17561 9180 17595
rect 9128 17552 9180 17561
rect 8300 17484 8352 17536
rect 8392 17484 8444 17536
rect 10692 17484 10744 17536
rect 12256 17595 12308 17604
rect 12256 17561 12265 17595
rect 12265 17561 12299 17595
rect 12299 17561 12308 17595
rect 12256 17552 12308 17561
rect 12716 17552 12768 17604
rect 16212 17552 16264 17604
rect 14096 17484 14148 17536
rect 14832 17527 14884 17536
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 14924 17484 14976 17536
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 20628 17620 20680 17672
rect 21180 17663 21232 17672
rect 21180 17629 21189 17663
rect 21189 17629 21223 17663
rect 21223 17629 21232 17663
rect 21180 17620 21232 17629
rect 22008 17620 22060 17672
rect 24032 17620 24084 17672
rect 29184 17688 29236 17740
rect 30196 17731 30248 17740
rect 30196 17697 30205 17731
rect 30205 17697 30239 17731
rect 30239 17697 30248 17731
rect 30196 17688 30248 17697
rect 30380 17756 30432 17808
rect 19616 17552 19668 17604
rect 18512 17484 18564 17536
rect 20444 17484 20496 17536
rect 20628 17484 20680 17536
rect 24400 17595 24452 17604
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 23572 17484 23624 17536
rect 24400 17561 24409 17595
rect 24409 17561 24443 17595
rect 24443 17561 24452 17595
rect 24400 17552 24452 17561
rect 25136 17595 25188 17604
rect 25136 17561 25145 17595
rect 25145 17561 25179 17595
rect 25179 17561 25188 17595
rect 25136 17552 25188 17561
rect 26792 17552 26844 17604
rect 27344 17595 27396 17604
rect 27344 17561 27353 17595
rect 27353 17561 27387 17595
rect 27387 17561 27396 17595
rect 27344 17552 27396 17561
rect 30840 17620 30892 17672
rect 31208 17620 31260 17672
rect 34704 17620 34756 17672
rect 30104 17595 30156 17604
rect 30104 17561 30113 17595
rect 30113 17561 30147 17595
rect 30147 17561 30156 17595
rect 30104 17552 30156 17561
rect 25228 17484 25280 17536
rect 27620 17484 27672 17536
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 28816 17484 28868 17493
rect 29184 17527 29236 17536
rect 29184 17493 29193 17527
rect 29193 17493 29227 17527
rect 29227 17493 29236 17527
rect 29184 17484 29236 17493
rect 30932 17527 30984 17536
rect 30932 17493 30941 17527
rect 30941 17493 30975 17527
rect 30975 17493 30984 17527
rect 30932 17484 30984 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 7380 17280 7432 17332
rect 8116 17280 8168 17332
rect 8392 17280 8444 17332
rect 9772 17280 9824 17332
rect 9864 17280 9916 17332
rect 12072 17280 12124 17332
rect 12532 17323 12584 17332
rect 12532 17289 12541 17323
rect 12541 17289 12575 17323
rect 12575 17289 12584 17323
rect 12532 17280 12584 17289
rect 14096 17280 14148 17332
rect 16120 17323 16172 17332
rect 16120 17289 16129 17323
rect 16129 17289 16163 17323
rect 16163 17289 16172 17323
rect 16120 17280 16172 17289
rect 17868 17280 17920 17332
rect 22836 17280 22888 17332
rect 23572 17280 23624 17332
rect 24216 17280 24268 17332
rect 4988 17212 5040 17264
rect 6460 17212 6512 17264
rect 12900 17255 12952 17264
rect 12900 17221 12909 17255
rect 12909 17221 12943 17255
rect 12943 17221 12952 17255
rect 12900 17212 12952 17221
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 1308 17076 1360 17128
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 6184 17144 6236 17196
rect 6368 17144 6420 17196
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 9036 17144 9088 17196
rect 9588 17144 9640 17196
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10876 17144 10928 17196
rect 11152 17144 11204 17196
rect 18696 17212 18748 17264
rect 20168 17255 20220 17264
rect 20168 17221 20177 17255
rect 20177 17221 20211 17255
rect 20211 17221 20220 17255
rect 20168 17212 20220 17221
rect 21916 17212 21968 17264
rect 28816 17280 28868 17332
rect 30104 17280 30156 17332
rect 30288 17280 30340 17332
rect 26792 17255 26844 17264
rect 26792 17221 26801 17255
rect 26801 17221 26835 17255
rect 26835 17221 26844 17255
rect 26792 17212 26844 17221
rect 30196 17212 30248 17264
rect 5816 17119 5868 17128
rect 5816 17085 5825 17119
rect 5825 17085 5859 17119
rect 5859 17085 5868 17119
rect 5816 17076 5868 17085
rect 5908 17076 5960 17128
rect 6736 17008 6788 17060
rect 7564 17076 7616 17128
rect 8760 17076 8812 17128
rect 8944 17076 8996 17128
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 17132 17144 17184 17196
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 21824 17144 21876 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 27804 17187 27856 17196
rect 27804 17153 27813 17187
rect 27813 17153 27847 17187
rect 27847 17153 27856 17187
rect 27804 17144 27856 17153
rect 29184 17144 29236 17196
rect 30104 17144 30156 17196
rect 30840 17187 30892 17196
rect 30840 17153 30849 17187
rect 30849 17153 30883 17187
rect 30883 17153 30892 17187
rect 30840 17144 30892 17153
rect 4344 16940 4396 16992
rect 6184 16940 6236 16992
rect 7472 16940 7524 16992
rect 7564 16940 7616 16992
rect 7840 16940 7892 16992
rect 8760 16940 8812 16992
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 9772 17008 9824 17060
rect 13360 17076 13412 17128
rect 15476 17076 15528 17128
rect 15844 17076 15896 17128
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 10324 17008 10376 17060
rect 11796 17008 11848 17060
rect 12072 16940 12124 16992
rect 12440 16940 12492 16992
rect 12532 16940 12584 16992
rect 13268 16940 13320 16992
rect 15016 17008 15068 17060
rect 17040 17008 17092 17060
rect 18512 17076 18564 17128
rect 18788 17076 18840 17128
rect 20996 17076 21048 17128
rect 21088 17076 21140 17128
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 16948 16940 17000 16992
rect 20628 17008 20680 17060
rect 20720 17051 20772 17060
rect 20720 17017 20729 17051
rect 20729 17017 20763 17051
rect 20763 17017 20772 17051
rect 20720 17008 20772 17017
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 22652 17008 22704 17060
rect 24584 17076 24636 17128
rect 27712 17076 27764 17128
rect 30380 17076 30432 17128
rect 45284 17008 45336 17060
rect 20076 16940 20128 16992
rect 21088 16940 21140 16992
rect 21364 16940 21416 16992
rect 22744 16940 22796 16992
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 26148 16940 26200 16992
rect 27252 16940 27304 16992
rect 30104 16940 30156 16992
rect 30288 16940 30340 16992
rect 48780 16940 48832 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 5724 16736 5776 16788
rect 6184 16736 6236 16788
rect 7564 16736 7616 16788
rect 8024 16736 8076 16788
rect 10416 16668 10468 16720
rect 12256 16668 12308 16720
rect 12900 16668 12952 16720
rect 6736 16600 6788 16652
rect 1308 16464 1360 16516
rect 7656 16532 7708 16584
rect 8116 16532 8168 16584
rect 10140 16532 10192 16584
rect 11336 16600 11388 16652
rect 14372 16736 14424 16788
rect 18880 16736 18932 16788
rect 21180 16736 21232 16788
rect 30932 16736 30984 16788
rect 18512 16668 18564 16720
rect 15200 16600 15252 16652
rect 16304 16600 16356 16652
rect 17224 16600 17276 16652
rect 20352 16600 20404 16652
rect 20720 16600 20772 16652
rect 23572 16668 23624 16720
rect 25136 16668 25188 16720
rect 22836 16600 22888 16652
rect 23848 16600 23900 16652
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 25320 16600 25372 16652
rect 25872 16600 25924 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27252 16643 27304 16652
rect 27252 16609 27261 16643
rect 27261 16609 27295 16643
rect 27295 16609 27304 16643
rect 27252 16600 27304 16609
rect 28632 16668 28684 16720
rect 30840 16668 30892 16720
rect 31300 16600 31352 16652
rect 12348 16532 12400 16584
rect 12440 16532 12492 16584
rect 14832 16532 14884 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 16580 16532 16632 16584
rect 17316 16532 17368 16584
rect 5172 16507 5224 16516
rect 5172 16473 5181 16507
rect 5181 16473 5215 16507
rect 5215 16473 5224 16507
rect 5172 16464 5224 16473
rect 7748 16464 7800 16516
rect 6736 16396 6788 16448
rect 6920 16396 6972 16448
rect 9036 16464 9088 16516
rect 12164 16464 12216 16516
rect 12808 16464 12860 16516
rect 8760 16396 8812 16448
rect 9772 16396 9824 16448
rect 10416 16396 10468 16448
rect 11244 16439 11296 16448
rect 11244 16405 11253 16439
rect 11253 16405 11287 16439
rect 11287 16405 11296 16439
rect 11244 16396 11296 16405
rect 11704 16396 11756 16448
rect 15568 16464 15620 16516
rect 18328 16532 18380 16584
rect 18604 16532 18656 16584
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 21824 16532 21876 16584
rect 23296 16532 23348 16584
rect 24032 16532 24084 16584
rect 25044 16532 25096 16584
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 16488 16396 16540 16448
rect 16672 16396 16724 16448
rect 19524 16396 19576 16448
rect 21456 16507 21508 16516
rect 21456 16473 21465 16507
rect 21465 16473 21499 16507
rect 21499 16473 21508 16507
rect 21456 16464 21508 16473
rect 23848 16464 23900 16516
rect 24124 16464 24176 16516
rect 21640 16396 21692 16448
rect 22468 16396 22520 16448
rect 23480 16396 23532 16448
rect 23756 16396 23808 16448
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25044 16396 25096 16405
rect 25320 16396 25372 16448
rect 25412 16396 25464 16448
rect 27712 16532 27764 16584
rect 28632 16532 28684 16584
rect 28448 16464 28500 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 4896 16192 4948 16244
rect 7380 16192 7432 16244
rect 10140 16192 10192 16244
rect 10232 16235 10284 16244
rect 10232 16201 10241 16235
rect 10241 16201 10275 16235
rect 10275 16201 10284 16235
rect 10232 16192 10284 16201
rect 12440 16192 12492 16244
rect 21456 16192 21508 16244
rect 24032 16192 24084 16244
rect 24492 16235 24544 16244
rect 24492 16201 24501 16235
rect 24501 16201 24535 16235
rect 24535 16201 24544 16235
rect 24492 16192 24544 16201
rect 24952 16192 25004 16244
rect 26792 16192 26844 16244
rect 27620 16192 27672 16244
rect 28632 16192 28684 16244
rect 3332 16124 3384 16176
rect 5816 16124 5868 16176
rect 10600 16167 10652 16176
rect 10600 16133 10609 16167
rect 10609 16133 10643 16167
rect 10643 16133 10652 16167
rect 10600 16124 10652 16133
rect 12256 16167 12308 16176
rect 12256 16133 12265 16167
rect 12265 16133 12299 16167
rect 12299 16133 12308 16167
rect 12256 16124 12308 16133
rect 12716 16124 12768 16176
rect 1308 15988 1360 16040
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 3792 16056 3844 16108
rect 4068 15988 4120 16040
rect 5724 16031 5776 16040
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 7380 16056 7432 16108
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 8300 16056 8352 16108
rect 8484 16099 8536 16108
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 6184 15988 6236 16040
rect 6552 15988 6604 16040
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 7472 15988 7524 16040
rect 8208 15988 8260 16040
rect 9956 15988 10008 16040
rect 10416 15988 10468 16040
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 10324 15920 10376 15972
rect 10876 15920 10928 15972
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 13636 15920 13688 15972
rect 15108 15988 15160 16040
rect 17592 16056 17644 16108
rect 15292 15920 15344 15972
rect 15936 15920 15988 15972
rect 5632 15852 5684 15904
rect 8576 15852 8628 15904
rect 12072 15852 12124 15904
rect 12900 15852 12952 15904
rect 13912 15852 13964 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16856 15988 16908 16040
rect 17868 16099 17920 16108
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 17868 16056 17920 16065
rect 19156 16056 19208 16108
rect 20444 16167 20496 16176
rect 20444 16133 20453 16167
rect 20453 16133 20487 16167
rect 20487 16133 20496 16167
rect 20444 16124 20496 16133
rect 17316 15920 17368 15972
rect 17500 15920 17552 15972
rect 18880 16031 18932 16040
rect 18880 15997 18889 16031
rect 18889 15997 18923 16031
rect 18923 15997 18932 16031
rect 18880 15988 18932 15997
rect 21824 16124 21876 16176
rect 23480 16124 23532 16176
rect 24400 16167 24452 16176
rect 24400 16133 24409 16167
rect 24409 16133 24443 16167
rect 24443 16133 24452 16167
rect 24400 16124 24452 16133
rect 25044 16124 25096 16176
rect 25412 16124 25464 16176
rect 22928 16056 22980 16108
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 21364 15920 21416 15972
rect 21732 15988 21784 16040
rect 24032 15988 24084 16040
rect 25136 16031 25188 16040
rect 25136 15997 25145 16031
rect 25145 15997 25179 16031
rect 25179 15997 25188 16031
rect 25136 15988 25188 15997
rect 27252 15988 27304 16040
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 17132 15852 17184 15904
rect 18604 15852 18656 15904
rect 19616 15852 19668 15904
rect 20812 15852 20864 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 21548 15852 21600 15904
rect 23848 15920 23900 15972
rect 24308 15852 24360 15904
rect 29736 15920 29788 15972
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 7196 15648 7248 15700
rect 8668 15648 8720 15700
rect 10968 15648 11020 15700
rect 12808 15648 12860 15700
rect 13360 15648 13412 15700
rect 1308 15512 1360 15564
rect 6184 15580 6236 15632
rect 5540 15512 5592 15564
rect 3424 15444 3476 15496
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 6920 15512 6972 15521
rect 7196 15444 7248 15496
rect 7564 15580 7616 15632
rect 8300 15512 8352 15564
rect 9220 15512 9272 15564
rect 10876 15512 10928 15564
rect 12072 15623 12124 15632
rect 12072 15589 12081 15623
rect 12081 15589 12115 15623
rect 12115 15589 12124 15623
rect 12072 15580 12124 15589
rect 12164 15580 12216 15632
rect 8668 15444 8720 15496
rect 12900 15512 12952 15564
rect 13636 15444 13688 15496
rect 23940 15648 23992 15700
rect 24492 15691 24544 15700
rect 24492 15657 24501 15691
rect 24501 15657 24535 15691
rect 24535 15657 24544 15691
rect 24492 15648 24544 15657
rect 13820 15580 13872 15632
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15108 15444 15160 15496
rect 7564 15376 7616 15428
rect 9220 15419 9272 15428
rect 9220 15385 9229 15419
rect 9229 15385 9263 15419
rect 9263 15385 9272 15419
rect 9220 15376 9272 15385
rect 9864 15376 9916 15428
rect 9956 15419 10008 15428
rect 9956 15385 9965 15419
rect 9965 15385 9999 15419
rect 9999 15385 10008 15419
rect 9956 15376 10008 15385
rect 10968 15376 11020 15428
rect 11060 15376 11112 15428
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 4804 15308 4856 15360
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 7840 15308 7892 15360
rect 8668 15308 8720 15360
rect 10416 15308 10468 15360
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 11796 15308 11848 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 13268 15376 13320 15428
rect 17040 15555 17092 15564
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 19432 15512 19484 15564
rect 20628 15512 20680 15564
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 21732 15580 21784 15632
rect 21916 15580 21968 15632
rect 22100 15580 22152 15632
rect 17316 15419 17368 15428
rect 17316 15385 17325 15419
rect 17325 15385 17359 15419
rect 17359 15385 17368 15419
rect 17316 15376 17368 15385
rect 17776 15376 17828 15428
rect 18604 15376 18656 15428
rect 13360 15308 13412 15360
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 14556 15308 14608 15360
rect 15384 15308 15436 15360
rect 16580 15308 16632 15360
rect 17408 15308 17460 15360
rect 19892 15376 19944 15428
rect 19708 15308 19760 15360
rect 20444 15308 20496 15360
rect 21916 15444 21968 15496
rect 21916 15308 21968 15360
rect 24308 15512 24360 15564
rect 25228 15512 25280 15564
rect 23296 15444 23348 15496
rect 26056 15444 26108 15496
rect 23572 15376 23624 15428
rect 23940 15419 23992 15428
rect 23940 15385 23949 15419
rect 23949 15385 23983 15419
rect 23983 15385 23992 15419
rect 23940 15376 23992 15385
rect 26148 15376 26200 15428
rect 22744 15308 22796 15360
rect 23848 15308 23900 15360
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 26056 15308 26108 15360
rect 48688 15376 48740 15428
rect 49240 15308 49292 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 3516 15147 3568 15156
rect 3516 15113 3525 15147
rect 3525 15113 3559 15147
rect 3559 15113 3568 15147
rect 3516 15104 3568 15113
rect 4068 15104 4120 15156
rect 6920 15104 6972 15156
rect 8668 15104 8720 15156
rect 11244 15104 11296 15156
rect 12624 15104 12676 15156
rect 13084 15104 13136 15156
rect 16672 15104 16724 15156
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 22100 15104 22152 15156
rect 23572 15104 23624 15156
rect 23848 15104 23900 15156
rect 24952 15104 25004 15156
rect 26792 15104 26844 15156
rect 4712 15036 4764 15088
rect 6276 15036 6328 15088
rect 7748 15036 7800 15088
rect 8576 15079 8628 15088
rect 8576 15045 8585 15079
rect 8585 15045 8619 15079
rect 8619 15045 8628 15079
rect 8576 15036 8628 15045
rect 8852 15036 8904 15088
rect 9036 15036 9088 15088
rect 9864 15036 9916 15088
rect 10784 15079 10836 15088
rect 10784 15045 10793 15079
rect 10793 15045 10827 15079
rect 10827 15045 10836 15079
rect 10784 15036 10836 15045
rect 1308 14900 1360 14952
rect 4068 14968 4120 15020
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 5816 14968 5868 15020
rect 6184 14968 6236 15020
rect 9956 14968 10008 15020
rect 13268 15036 13320 15088
rect 14740 15036 14792 15088
rect 15108 15036 15160 15088
rect 15292 15036 15344 15088
rect 16580 15036 16632 15088
rect 19524 15036 19576 15088
rect 21640 15036 21692 15088
rect 22744 15036 22796 15088
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 12072 14968 12124 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 17592 14968 17644 15020
rect 19708 14968 19760 15020
rect 19984 14968 20036 15020
rect 7288 14900 7340 14952
rect 7656 14900 7708 14952
rect 3608 14832 3660 14884
rect 4068 14832 4120 14884
rect 4436 14764 4488 14816
rect 6828 14764 6880 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 8300 14832 8352 14884
rect 9496 14832 9548 14884
rect 11336 14900 11388 14952
rect 12256 14900 12308 14952
rect 14280 14900 14332 14952
rect 10048 14764 10100 14816
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 13728 14832 13780 14884
rect 16120 14900 16172 14952
rect 19248 14900 19300 14952
rect 15844 14832 15896 14884
rect 17592 14832 17644 14884
rect 17868 14832 17920 14884
rect 19616 14832 19668 14884
rect 19708 14875 19760 14884
rect 19708 14841 19717 14875
rect 19717 14841 19751 14875
rect 19751 14841 19760 14875
rect 19708 14832 19760 14841
rect 20628 14968 20680 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23940 14968 23992 15020
rect 22652 14900 22704 14952
rect 21916 14832 21968 14884
rect 14188 14764 14240 14816
rect 15292 14764 15344 14816
rect 16304 14807 16356 14816
rect 16304 14773 16313 14807
rect 16313 14773 16347 14807
rect 16347 14773 16356 14807
rect 16304 14764 16356 14773
rect 17776 14764 17828 14816
rect 18880 14764 18932 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 19524 14764 19576 14816
rect 24860 14832 24912 14884
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 4160 14560 4212 14612
rect 4712 14560 4764 14612
rect 4896 14560 4948 14612
rect 4988 14560 5040 14612
rect 9220 14560 9272 14612
rect 10692 14560 10744 14612
rect 10784 14560 10836 14612
rect 7196 14535 7248 14544
rect 7196 14501 7205 14535
rect 7205 14501 7239 14535
rect 7239 14501 7248 14535
rect 7196 14492 7248 14501
rect 7656 14492 7708 14544
rect 1308 14424 1360 14476
rect 4252 14424 4304 14476
rect 4436 14424 4488 14476
rect 6736 14424 6788 14476
rect 9864 14492 9916 14544
rect 10048 14492 10100 14544
rect 10140 14492 10192 14544
rect 5172 14356 5224 14408
rect 7196 14356 7248 14408
rect 7840 14356 7892 14408
rect 8668 14424 8720 14476
rect 9680 14424 9732 14476
rect 10232 14424 10284 14476
rect 9772 14356 9824 14408
rect 10876 14356 10928 14408
rect 11060 14356 11112 14408
rect 4160 14220 4212 14272
rect 5816 14288 5868 14340
rect 6276 14288 6328 14340
rect 9404 14288 9456 14340
rect 9680 14288 9732 14340
rect 10140 14288 10192 14340
rect 10232 14288 10284 14340
rect 13544 14560 13596 14612
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 14464 14560 14516 14612
rect 15108 14560 15160 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 21088 14560 21140 14612
rect 34888 14560 34940 14612
rect 12256 14424 12308 14476
rect 12808 14424 12860 14476
rect 12900 14424 12952 14476
rect 14188 14424 14240 14476
rect 16304 14424 16356 14476
rect 17132 14424 17184 14476
rect 17224 14424 17276 14476
rect 18328 14424 18380 14476
rect 19248 14424 19300 14476
rect 22008 14424 22060 14476
rect 23940 14424 23992 14476
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 14280 14356 14332 14408
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8760 14220 8812 14272
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 9864 14220 9916 14272
rect 12256 14331 12308 14340
rect 12256 14297 12265 14331
rect 12265 14297 12299 14331
rect 12299 14297 12308 14331
rect 12256 14288 12308 14297
rect 12716 14288 12768 14340
rect 13176 14220 13228 14272
rect 15384 14288 15436 14340
rect 16856 14288 16908 14340
rect 17408 14288 17460 14340
rect 17868 14288 17920 14340
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 16488 14220 16540 14272
rect 26608 14424 26660 14476
rect 21088 14288 21140 14340
rect 21916 14288 21968 14340
rect 23848 14288 23900 14340
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 21456 14220 21508 14272
rect 21824 14220 21876 14272
rect 22744 14220 22796 14272
rect 26148 14399 26200 14408
rect 26148 14365 26157 14399
rect 26157 14365 26191 14399
rect 26191 14365 26200 14399
rect 26148 14356 26200 14365
rect 24952 14331 25004 14340
rect 24952 14297 24961 14331
rect 24961 14297 24995 14331
rect 24995 14297 25004 14331
rect 24952 14288 25004 14297
rect 25044 14331 25096 14340
rect 25044 14297 25053 14331
rect 25053 14297 25087 14331
rect 25087 14297 25096 14331
rect 25044 14288 25096 14297
rect 25320 14288 25372 14340
rect 24308 14220 24360 14272
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 25688 14220 25740 14272
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 26148 14220 26200 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 4160 14016 4212 14068
rect 4988 14016 5040 14068
rect 6368 14016 6420 14068
rect 4252 13948 4304 14000
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7380 14059 7432 14068
rect 7380 14025 7389 14059
rect 7389 14025 7423 14059
rect 7423 14025 7432 14059
rect 7380 14016 7432 14025
rect 9220 14016 9272 14068
rect 11428 14016 11480 14068
rect 8576 13991 8628 14000
rect 8576 13957 8585 13991
rect 8585 13957 8619 13991
rect 8619 13957 8628 13991
rect 8576 13948 8628 13957
rect 10600 13948 10652 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 5632 13880 5684 13932
rect 6276 13880 6328 13932
rect 1308 13812 1360 13864
rect 2504 13812 2556 13864
rect 4896 13812 4948 13864
rect 5448 13812 5500 13864
rect 7288 13812 7340 13864
rect 7656 13880 7708 13932
rect 11704 14016 11756 14068
rect 12072 14016 12124 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 13544 14016 13596 14068
rect 17224 14016 17276 14068
rect 17316 14016 17368 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 19616 14016 19668 14068
rect 21180 14016 21232 14068
rect 25780 14016 25832 14068
rect 11796 13948 11848 14000
rect 12072 13880 12124 13932
rect 12348 13880 12400 13932
rect 5908 13744 5960 13796
rect 7656 13744 7708 13796
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 10048 13812 10100 13864
rect 11520 13812 11572 13864
rect 11796 13812 11848 13864
rect 12164 13812 12216 13864
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 16672 13948 16724 14000
rect 17868 13948 17920 14000
rect 20996 13948 21048 14000
rect 12808 13812 12860 13864
rect 15200 13880 15252 13932
rect 16948 13880 17000 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 10600 13744 10652 13796
rect 13636 13744 13688 13796
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 5448 13676 5500 13728
rect 5816 13676 5868 13728
rect 7472 13676 7524 13728
rect 8944 13676 8996 13728
rect 9036 13676 9088 13728
rect 9404 13676 9456 13728
rect 12348 13676 12400 13728
rect 14464 13744 14516 13796
rect 15108 13812 15160 13864
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 17776 13812 17828 13864
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 21640 13880 21692 13932
rect 21824 13948 21876 14000
rect 22008 13880 22060 13932
rect 24584 13948 24636 14000
rect 25320 13948 25372 14000
rect 25688 13948 25740 14000
rect 16304 13676 16356 13728
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 20720 13744 20772 13796
rect 18972 13676 19024 13728
rect 20168 13676 20220 13728
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 24124 13744 24176 13796
rect 21916 13676 21968 13728
rect 22560 13676 22612 13728
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 5172 13472 5224 13524
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 5172 13336 5224 13388
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 7748 13472 7800 13524
rect 10140 13472 10192 13524
rect 10692 13472 10744 13524
rect 7380 13336 7432 13388
rect 7748 13336 7800 13388
rect 9036 13336 9088 13388
rect 10600 13404 10652 13456
rect 11060 13404 11112 13456
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 6276 13268 6328 13320
rect 3332 13243 3384 13252
rect 3332 13209 3341 13243
rect 3341 13209 3375 13243
rect 3375 13209 3384 13243
rect 3332 13200 3384 13209
rect 4436 13243 4488 13252
rect 4436 13209 4445 13243
rect 4445 13209 4479 13243
rect 4479 13209 4488 13243
rect 4436 13200 4488 13209
rect 1860 13132 1912 13184
rect 6920 13200 6972 13252
rect 7288 13200 7340 13252
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6276 13132 6328 13184
rect 7656 13132 7708 13184
rect 8760 13200 8812 13252
rect 9588 13200 9640 13252
rect 9680 13200 9732 13252
rect 9496 13132 9548 13184
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 12256 13472 12308 13524
rect 15016 13472 15068 13524
rect 17408 13472 17460 13524
rect 18788 13404 18840 13456
rect 21916 13472 21968 13524
rect 22652 13472 22704 13524
rect 23112 13472 23164 13524
rect 24492 13472 24544 13524
rect 21640 13404 21692 13456
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 13268 13336 13320 13388
rect 15200 13336 15252 13388
rect 16396 13336 16448 13388
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 17868 13336 17920 13388
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 12256 13243 12308 13252
rect 12256 13209 12265 13243
rect 12265 13209 12299 13243
rect 12299 13209 12308 13243
rect 12256 13200 12308 13209
rect 12716 13200 12768 13252
rect 14188 13200 14240 13252
rect 16304 13200 16356 13252
rect 14648 13132 14700 13184
rect 17868 13200 17920 13252
rect 18328 13132 18380 13184
rect 22192 13336 22244 13388
rect 23756 13404 23808 13456
rect 23848 13404 23900 13456
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 23572 13336 23624 13388
rect 32496 13336 32548 13388
rect 21732 13268 21784 13320
rect 22008 13268 22060 13320
rect 23020 13268 23072 13320
rect 18972 13200 19024 13252
rect 20352 13132 20404 13184
rect 22928 13132 22980 13184
rect 24492 13200 24544 13252
rect 29736 13200 29788 13252
rect 25228 13132 25280 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6552 12928 6604 12980
rect 7104 12928 7156 12980
rect 9864 12928 9916 12980
rect 10140 12928 10192 12980
rect 10692 12928 10744 12980
rect 11152 12928 11204 12980
rect 3700 12903 3752 12912
rect 3700 12869 3709 12903
rect 3709 12869 3743 12903
rect 3743 12869 3752 12903
rect 3700 12860 3752 12869
rect 4344 12860 4396 12912
rect 5816 12860 5868 12912
rect 7012 12860 7064 12912
rect 8576 12860 8628 12912
rect 8760 12860 8812 12912
rect 9588 12860 9640 12912
rect 12440 12860 12492 12912
rect 1308 12792 1360 12844
rect 3792 12792 3844 12844
rect 4436 12792 4488 12844
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 3424 12724 3476 12776
rect 3700 12724 3752 12776
rect 6920 12792 6972 12844
rect 10324 12792 10376 12844
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 7748 12656 7800 12708
rect 5632 12588 5684 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7380 12588 7432 12640
rect 9036 12724 9088 12776
rect 10140 12724 10192 12776
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 15384 12928 15436 12980
rect 16948 12928 17000 12980
rect 20168 12928 20220 12980
rect 21180 12928 21232 12980
rect 21732 12928 21784 12980
rect 22928 12928 22980 12980
rect 23480 12928 23532 12980
rect 13268 12792 13320 12844
rect 14280 12860 14332 12912
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 18420 12860 18472 12912
rect 18880 12860 18932 12912
rect 19156 12860 19208 12912
rect 23572 12860 23624 12912
rect 23940 12860 23992 12912
rect 14924 12792 14976 12801
rect 18696 12792 18748 12844
rect 21548 12792 21600 12844
rect 22192 12792 22244 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 14280 12724 14332 12776
rect 15108 12724 15160 12776
rect 15200 12724 15252 12776
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 14924 12656 14976 12708
rect 18512 12656 18564 12708
rect 20076 12724 20128 12776
rect 21456 12724 21508 12776
rect 24308 12724 24360 12776
rect 9312 12588 9364 12640
rect 11612 12631 11664 12640
rect 11612 12597 11621 12631
rect 11621 12597 11655 12631
rect 11655 12597 11664 12631
rect 11612 12588 11664 12597
rect 12164 12588 12216 12640
rect 13268 12588 13320 12640
rect 14556 12588 14608 12640
rect 15292 12588 15344 12640
rect 16672 12588 16724 12640
rect 17040 12588 17092 12640
rect 18696 12588 18748 12640
rect 22468 12656 22520 12708
rect 20904 12588 20956 12640
rect 23940 12588 23992 12640
rect 24400 12588 24452 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 2872 12384 2924 12436
rect 4344 12384 4396 12436
rect 4712 12384 4764 12436
rect 9680 12384 9732 12436
rect 4528 12248 4580 12300
rect 7288 12316 7340 12368
rect 5172 12248 5224 12300
rect 7748 12248 7800 12300
rect 8208 12316 8260 12368
rect 9312 12248 9364 12300
rect 1308 12180 1360 12232
rect 4160 12223 4212 12232
rect 1952 12112 2004 12164
rect 2504 12112 2556 12164
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 4344 12180 4396 12232
rect 4804 12180 4856 12232
rect 7472 12180 7524 12232
rect 8208 12180 8260 12232
rect 10416 12180 10468 12232
rect 11612 12316 11664 12368
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 12532 12384 12584 12436
rect 14188 12427 14240 12436
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 14280 12384 14332 12436
rect 14096 12316 14148 12368
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 18788 12384 18840 12436
rect 20720 12384 20772 12436
rect 11796 12248 11848 12300
rect 12256 12248 12308 12300
rect 19892 12316 19944 12368
rect 15200 12248 15252 12300
rect 15384 12248 15436 12300
rect 16212 12248 16264 12300
rect 17040 12248 17092 12300
rect 18328 12291 18380 12300
rect 18328 12257 18337 12291
rect 18337 12257 18371 12291
rect 18371 12257 18380 12291
rect 18328 12248 18380 12257
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 20352 12291 20404 12300
rect 20352 12257 20361 12291
rect 20361 12257 20395 12291
rect 20395 12257 20404 12291
rect 20352 12248 20404 12257
rect 24400 12427 24452 12436
rect 24400 12393 24409 12427
rect 24409 12393 24443 12427
rect 24443 12393 24452 12427
rect 24400 12384 24452 12393
rect 14924 12180 14976 12232
rect 5540 12112 5592 12164
rect 5724 12112 5776 12164
rect 6276 12112 6328 12164
rect 9128 12155 9180 12164
rect 9128 12121 9137 12155
rect 9137 12121 9171 12155
rect 9171 12121 9180 12155
rect 9128 12112 9180 12121
rect 9956 12112 10008 12164
rect 6920 12044 6972 12096
rect 8944 12044 8996 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10692 12044 10744 12096
rect 11244 12044 11296 12096
rect 12072 12044 12124 12096
rect 12256 12087 12308 12096
rect 12256 12053 12265 12087
rect 12265 12053 12299 12087
rect 12299 12053 12308 12087
rect 12256 12044 12308 12053
rect 13268 12044 13320 12096
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 14464 12112 14516 12164
rect 17040 12112 17092 12164
rect 17408 12044 17460 12096
rect 18328 12112 18380 12164
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 18880 12155 18932 12164
rect 18880 12121 18889 12155
rect 18889 12121 18923 12155
rect 18923 12121 18932 12155
rect 18880 12112 18932 12121
rect 19248 12044 19300 12096
rect 22192 12180 22244 12232
rect 23940 12180 23992 12232
rect 21732 12112 21784 12164
rect 25044 12112 25096 12164
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 1308 11840 1360 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 2320 11704 2372 11756
rect 5264 11704 5316 11756
rect 6828 11772 6880 11824
rect 7656 11815 7708 11824
rect 7656 11781 7665 11815
rect 7665 11781 7699 11815
rect 7699 11781 7708 11815
rect 7656 11772 7708 11781
rect 8208 11772 8260 11824
rect 6552 11704 6604 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 9956 11704 10008 11756
rect 12256 11840 12308 11892
rect 12808 11840 12860 11892
rect 15200 11883 15252 11892
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 10600 11772 10652 11824
rect 13360 11772 13412 11824
rect 14188 11772 14240 11824
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 17776 11840 17828 11892
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 14740 11704 14792 11756
rect 16120 11704 16172 11756
rect 17592 11772 17644 11824
rect 20904 11840 20956 11892
rect 21732 11840 21784 11892
rect 1952 11636 2004 11688
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 2780 11636 2832 11688
rect 4068 11636 4120 11688
rect 5632 11636 5684 11688
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 7196 11636 7248 11688
rect 8116 11636 8168 11688
rect 5540 11568 5592 11620
rect 7012 11568 7064 11620
rect 7380 11568 7432 11620
rect 7656 11500 7708 11552
rect 7840 11500 7892 11552
rect 9036 11568 9088 11620
rect 11796 11636 11848 11688
rect 12256 11636 12308 11688
rect 15016 11636 15068 11688
rect 17040 11636 17092 11688
rect 11520 11568 11572 11620
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 8760 11500 8812 11552
rect 10508 11500 10560 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12072 11500 12124 11552
rect 15016 11500 15068 11552
rect 15292 11500 15344 11552
rect 18512 11568 18564 11620
rect 19708 11679 19760 11688
rect 19708 11645 19717 11679
rect 19717 11645 19751 11679
rect 19751 11645 19760 11679
rect 19708 11636 19760 11645
rect 24032 11840 24084 11892
rect 24400 11883 24452 11892
rect 24400 11849 24409 11883
rect 24409 11849 24443 11883
rect 24443 11849 24452 11883
rect 24400 11840 24452 11849
rect 22744 11772 22796 11824
rect 23940 11772 23992 11824
rect 22192 11636 22244 11688
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 2780 11228 2832 11280
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 3424 11296 3476 11348
rect 3608 11296 3660 11348
rect 5540 11296 5592 11348
rect 5724 11296 5776 11348
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 3608 11203 3660 11212
rect 3608 11169 3617 11203
rect 3617 11169 3651 11203
rect 3651 11169 3660 11203
rect 3608 11160 3660 11169
rect 6828 11160 6880 11212
rect 6368 11092 6420 11144
rect 6736 11092 6788 11144
rect 12532 11296 12584 11348
rect 13452 11296 13504 11348
rect 14188 11296 14240 11348
rect 7748 11228 7800 11280
rect 8760 11228 8812 11280
rect 9036 11228 9088 11280
rect 8116 11160 8168 11212
rect 9220 11160 9272 11212
rect 12808 11228 12860 11280
rect 16120 11296 16172 11348
rect 16212 11296 16264 11348
rect 18972 11296 19024 11348
rect 22836 11296 22888 11348
rect 23940 11296 23992 11348
rect 30104 11296 30156 11348
rect 9772 11160 9824 11212
rect 10232 11160 10284 11212
rect 8300 11092 8352 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 7932 11024 7984 11076
rect 6736 10956 6788 11008
rect 8208 10956 8260 11008
rect 9404 11024 9456 11076
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 12348 11160 12400 11212
rect 13360 11160 13412 11212
rect 19984 11160 20036 11212
rect 29736 11203 29788 11212
rect 29736 11169 29745 11203
rect 29745 11169 29779 11203
rect 29779 11169 29788 11203
rect 29736 11160 29788 11169
rect 14464 11092 14516 11144
rect 16856 11092 16908 11144
rect 19248 11092 19300 11144
rect 9220 10956 9272 11008
rect 10324 10999 10376 11008
rect 10324 10965 10333 10999
rect 10333 10965 10367 10999
rect 10367 10965 10376 10999
rect 10324 10956 10376 10965
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 13452 11024 13504 11076
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 17316 11024 17368 11076
rect 12440 10956 12492 11008
rect 15200 10956 15252 11008
rect 17868 11024 17920 11076
rect 19708 11024 19760 11076
rect 31300 11092 31352 11144
rect 47860 11092 47912 11144
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 21732 11024 21784 11076
rect 27804 11024 27856 11076
rect 30104 11024 30156 11076
rect 17776 10956 17828 11008
rect 18420 10956 18472 11008
rect 20628 10956 20680 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 3608 10752 3660 10804
rect 6736 10684 6788 10736
rect 8300 10684 8352 10736
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 10968 10752 11020 10804
rect 11520 10752 11572 10804
rect 12256 10752 12308 10804
rect 12072 10684 12124 10736
rect 15292 10752 15344 10804
rect 17040 10752 17092 10804
rect 15660 10684 15712 10736
rect 15752 10684 15804 10736
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 5264 10616 5316 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 13452 10616 13504 10668
rect 4988 10548 5040 10600
rect 7380 10548 7432 10600
rect 7012 10480 7064 10532
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 7380 10412 7432 10464
rect 8116 10548 8168 10600
rect 8760 10548 8812 10600
rect 10048 10548 10100 10600
rect 11244 10548 11296 10600
rect 12348 10548 12400 10600
rect 15384 10616 15436 10668
rect 15200 10548 15252 10600
rect 7840 10412 7892 10464
rect 8208 10412 8260 10464
rect 14832 10480 14884 10532
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 16304 10548 16356 10600
rect 17868 10684 17920 10736
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 21456 10752 21508 10804
rect 21732 10752 21784 10804
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 22836 10548 22888 10600
rect 9036 10412 9088 10464
rect 9496 10412 9548 10464
rect 10508 10412 10560 10464
rect 14004 10412 14056 10464
rect 20536 10412 20588 10464
rect 20628 10412 20680 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 3792 10208 3844 10260
rect 6736 10208 6788 10260
rect 7564 10208 7616 10260
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 10784 10208 10836 10260
rect 10968 10208 11020 10260
rect 22284 10208 22336 10260
rect 8116 10140 8168 10192
rect 10876 10140 10928 10192
rect 13452 10140 13504 10192
rect 13820 10140 13872 10192
rect 1584 10115 1636 10124
rect 1584 10081 1593 10115
rect 1593 10081 1627 10115
rect 1627 10081 1636 10115
rect 1584 10072 1636 10081
rect 3700 10072 3752 10124
rect 3884 10072 3936 10124
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 7840 10072 7892 10124
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 11980 10072 12032 10124
rect 4068 10004 4120 10056
rect 4436 10004 4488 10056
rect 3792 9936 3844 9988
rect 7196 9936 7248 9988
rect 7564 9936 7616 9988
rect 10968 9936 11020 9988
rect 9128 9868 9180 9920
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 11520 9979 11572 9988
rect 11520 9945 11529 9979
rect 11529 9945 11563 9979
rect 11563 9945 11572 9979
rect 11520 9936 11572 9945
rect 19156 10140 19208 10192
rect 15200 10072 15252 10124
rect 16212 10072 16264 10124
rect 14464 10004 14516 10056
rect 16856 10004 16908 10056
rect 19708 10072 19760 10124
rect 20168 10072 20220 10124
rect 21732 10140 21784 10192
rect 15292 9936 15344 9988
rect 17040 9936 17092 9988
rect 11796 9868 11848 9920
rect 11888 9868 11940 9920
rect 15016 9868 15068 9920
rect 16488 9868 16540 9920
rect 19708 9979 19760 9988
rect 19708 9945 19717 9979
rect 19717 9945 19751 9979
rect 19751 9945 19760 9979
rect 19708 9936 19760 9945
rect 18328 9868 18380 9920
rect 24124 9936 24176 9988
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1492 9707 1544 9716
rect 1492 9673 1501 9707
rect 1501 9673 1535 9707
rect 1535 9673 1544 9707
rect 1492 9664 1544 9673
rect 7380 9664 7432 9716
rect 13636 9664 13688 9716
rect 13820 9707 13872 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 6000 9596 6052 9648
rect 8668 9596 8720 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 13820 9673 13829 9707
rect 13829 9673 13863 9707
rect 13863 9673 13872 9707
rect 13820 9664 13872 9673
rect 16212 9707 16264 9716
rect 16212 9673 16221 9707
rect 16221 9673 16255 9707
rect 16255 9673 16264 9707
rect 16212 9664 16264 9673
rect 16488 9596 16540 9648
rect 18420 9664 18472 9716
rect 19156 9664 19208 9716
rect 18696 9596 18748 9648
rect 24584 9596 24636 9648
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 5172 9528 5224 9580
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 7840 9528 7892 9580
rect 9496 9528 9548 9580
rect 9680 9528 9732 9580
rect 1676 9460 1728 9512
rect 2596 9460 2648 9512
rect 4528 9503 4580 9512
rect 4528 9469 4537 9503
rect 4537 9469 4571 9503
rect 4571 9469 4580 9503
rect 4528 9460 4580 9469
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7748 9460 7800 9512
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11244 9460 11296 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 3608 9435 3660 9444
rect 3608 9401 3617 9435
rect 3617 9401 3651 9435
rect 3651 9401 3660 9435
rect 3608 9392 3660 9401
rect 13544 9392 13596 9444
rect 16672 9460 16724 9512
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17132 9460 17184 9512
rect 17224 9460 17276 9512
rect 27528 9571 27580 9580
rect 27528 9537 27537 9571
rect 27537 9537 27571 9571
rect 27571 9537 27580 9571
rect 27528 9528 27580 9537
rect 21180 9460 21232 9512
rect 22560 9460 22612 9512
rect 7196 9324 7248 9376
rect 8760 9324 8812 9376
rect 11612 9324 11664 9376
rect 12440 9324 12492 9376
rect 14556 9324 14608 9376
rect 18328 9392 18380 9444
rect 19064 9435 19116 9444
rect 19064 9401 19073 9435
rect 19073 9401 19107 9435
rect 19107 9401 19116 9435
rect 19064 9392 19116 9401
rect 16120 9324 16172 9376
rect 18696 9324 18748 9376
rect 20168 9324 20220 9376
rect 31300 9596 31352 9648
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 2688 9120 2740 9172
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 9680 9120 9732 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 32864 9120 32916 9172
rect 6828 9052 6880 9104
rect 2872 8916 2924 8968
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 5540 8916 5592 8968
rect 7748 8916 7800 8968
rect 7932 8916 7984 8968
rect 8668 9052 8720 9104
rect 10048 9052 10100 9104
rect 8760 8984 8812 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9588 8984 9640 9036
rect 11980 9052 12032 9104
rect 14740 9052 14792 9104
rect 10232 8916 10284 8968
rect 10324 8916 10376 8968
rect 11796 8984 11848 9036
rect 15476 9052 15528 9104
rect 15752 8984 15804 9036
rect 16856 8984 16908 9036
rect 9128 8848 9180 8900
rect 6644 8780 6696 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 9496 8848 9548 8900
rect 10048 8848 10100 8900
rect 11888 8848 11940 8900
rect 11980 8848 12032 8900
rect 13176 8848 13228 8900
rect 9680 8780 9732 8832
rect 12532 8780 12584 8832
rect 13360 8916 13412 8968
rect 16212 8848 16264 8900
rect 15016 8780 15068 8832
rect 16672 8780 16724 8832
rect 17592 8780 17644 8832
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 3332 8619 3384 8628
rect 3332 8585 3341 8619
rect 3341 8585 3375 8619
rect 3375 8585 3384 8619
rect 3332 8576 3384 8585
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 5264 8576 5316 8628
rect 7288 8619 7340 8628
rect 7288 8585 7297 8619
rect 7297 8585 7331 8619
rect 7331 8585 7340 8619
rect 7288 8576 7340 8585
rect 7380 8576 7432 8628
rect 9588 8576 9640 8628
rect 12348 8576 12400 8628
rect 12532 8619 12584 8628
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 15384 8576 15436 8628
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 5172 8508 5224 8517
rect 5356 8508 5408 8560
rect 11796 8508 11848 8560
rect 16304 8576 16356 8628
rect 20444 8508 20496 8560
rect 2780 8440 2832 8492
rect 3332 8440 3384 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4988 8440 5040 8492
rect 6368 8440 6420 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 6460 8372 6512 8424
rect 4344 8304 4396 8356
rect 8576 8440 8628 8492
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 6920 8304 6972 8356
rect 9588 8347 9640 8356
rect 9588 8313 9597 8347
rect 9597 8313 9631 8347
rect 9631 8313 9640 8347
rect 9588 8304 9640 8313
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 13544 8440 13596 8492
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 14556 8372 14608 8424
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 18420 8440 18472 8492
rect 11060 8304 11112 8356
rect 12440 8304 12492 8356
rect 20352 8372 20404 8424
rect 13360 8236 13412 8288
rect 14740 8236 14792 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1676 8032 1728 8084
rect 3424 8032 3476 8084
rect 4160 8032 4212 8084
rect 8300 8032 8352 8084
rect 9956 8032 10008 8084
rect 3700 7896 3752 7948
rect 2872 7828 2924 7880
rect 8392 7964 8444 8016
rect 11704 7964 11756 8016
rect 10140 7939 10192 7948
rect 10140 7905 10149 7939
rect 10149 7905 10183 7939
rect 10183 7905 10192 7939
rect 10140 7896 10192 7905
rect 11152 7896 11204 7948
rect 11336 7896 11388 7948
rect 17224 8032 17276 8084
rect 11980 7964 12032 8016
rect 13360 7896 13412 7948
rect 3424 7760 3476 7812
rect 11428 7828 11480 7880
rect 13728 7896 13780 7948
rect 15200 8007 15252 8016
rect 15200 7973 15209 8007
rect 15209 7973 15243 8007
rect 15243 7973 15252 8007
rect 15200 7964 15252 7973
rect 22560 7828 22612 7880
rect 6092 7692 6144 7744
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 19708 7760 19760 7812
rect 16580 7692 16632 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 1952 7488 2004 7540
rect 2044 7488 2096 7540
rect 1860 7352 1912 7404
rect 3332 7488 3384 7540
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 13360 7488 13412 7540
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 27804 7488 27856 7540
rect 9220 7420 9272 7472
rect 2504 7352 2556 7404
rect 2780 7284 2832 7336
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 11612 7420 11664 7472
rect 24032 7420 24084 7472
rect 3332 7284 3384 7336
rect 7656 7284 7708 7336
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22468 7327 22520 7336
rect 22468 7293 22477 7327
rect 22477 7293 22511 7327
rect 22511 7293 22520 7327
rect 22468 7284 22520 7293
rect 15660 7216 15712 7268
rect 9036 7148 9088 7200
rect 14004 7148 14056 7200
rect 17500 7148 17552 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 2780 6876 2832 6928
rect 23940 6944 23992 6996
rect 8852 6808 8904 6860
rect 10508 6808 10560 6860
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 1308 6672 1360 6724
rect 20904 6740 20956 6792
rect 27528 6740 27580 6792
rect 1400 6604 1452 6656
rect 10692 6672 10744 6724
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 22100 6604 22152 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 1768 6400 1820 6452
rect 3976 6400 4028 6452
rect 2872 6264 2924 6316
rect 22560 6264 22612 6316
rect 1308 6196 1360 6248
rect 12164 6196 12216 6248
rect 7472 6128 7524 6180
rect 24860 6060 24912 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 1308 5856 1360 5908
rect 22468 5856 22520 5908
rect 12808 5788 12860 5840
rect 14004 5720 14056 5772
rect 16856 5720 16908 5772
rect 22100 5720 22152 5772
rect 24860 5763 24912 5772
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 28724 5720 28776 5772
rect 1308 5652 1360 5704
rect 9772 5652 9824 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 16580 5584 16632 5636
rect 18696 5584 18748 5636
rect 25504 5584 25556 5636
rect 17040 5516 17092 5568
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 27160 5627 27212 5636
rect 27160 5593 27169 5627
rect 27169 5593 27203 5627
rect 27203 5593 27212 5627
rect 27160 5584 27212 5593
rect 27344 5584 27396 5636
rect 27528 5584 27580 5636
rect 28908 5584 28960 5636
rect 27620 5516 27672 5568
rect 28540 5516 28592 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 27160 5312 27212 5364
rect 28356 5244 28408 5296
rect 1308 5176 1360 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 9864 5108 9916 5160
rect 15476 5108 15528 5160
rect 21364 5176 21416 5228
rect 22100 5219 22152 5228
rect 22100 5185 22144 5219
rect 22144 5185 22152 5219
rect 22100 5176 22152 5185
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 28816 5151 28868 5160
rect 28816 5117 28825 5151
rect 28825 5117 28859 5151
rect 28859 5117 28868 5151
rect 28816 5108 28868 5117
rect 41420 5108 41472 5160
rect 33508 5040 33560 5092
rect 17868 4972 17920 5024
rect 20536 4972 20588 5024
rect 25964 4972 26016 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 16580 4768 16632 4820
rect 28816 4768 28868 4820
rect 1308 4632 1360 4684
rect 11520 4632 11572 4684
rect 25964 4675 26016 4684
rect 25964 4641 25973 4675
rect 25973 4641 26007 4675
rect 26007 4641 26016 4675
rect 25964 4632 26016 4641
rect 27528 4675 27580 4684
rect 27528 4641 27537 4675
rect 27537 4641 27571 4675
rect 27571 4641 27580 4675
rect 27528 4632 27580 4641
rect 20904 4564 20956 4616
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 17684 4428 17736 4480
rect 27804 4428 27856 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 2780 4156 2832 4208
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2872 4088 2924 4140
rect 2688 3952 2740 4004
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 6276 4088 6328 4140
rect 10600 4088 10652 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 9956 3952 10008 4004
rect 9680 3884 9732 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 1308 3680 1360 3732
rect 2780 3680 2832 3732
rect 11428 3680 11480 3732
rect 1308 3476 1360 3528
rect 28908 3612 28960 3664
rect 44088 3612 44140 3664
rect 7012 3544 7064 3596
rect 27528 3544 27580 3596
rect 46756 3544 46808 3596
rect 11980 3476 12032 3528
rect 28540 3476 28592 3528
rect 49424 3476 49476 3528
rect 3424 3408 3476 3460
rect 12624 3408 12676 3460
rect 19340 3408 19392 3460
rect 38752 3408 38804 3460
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 3424 3136 3476 3188
rect 8300 3136 8352 3188
rect 6920 3068 6972 3120
rect 10048 3068 10100 3120
rect 12808 3068 12860 3120
rect 15476 3068 15528 3120
rect 17684 3068 17736 3120
rect 2780 3000 2832 3052
rect 7840 3000 7892 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17868 3000 17920 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 1308 2932 1360 2984
rect 7196 2932 7248 2984
rect 9772 2932 9824 2984
rect 1400 2796 1452 2848
rect 2872 2796 2924 2848
rect 10048 2796 10100 2848
rect 12440 2864 12492 2916
rect 16580 2796 16632 2848
rect 17500 2796 17552 2848
rect 20076 2796 20128 2848
rect 22008 2796 22060 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 7196 2592 7248 2644
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 27804 2592 27856 2644
rect 28724 2592 28776 2644
rect 33508 2635 33560 2644
rect 33508 2601 33517 2635
rect 33517 2601 33551 2635
rect 33551 2601 33560 2635
rect 33508 2592 33560 2601
rect 1308 2456 1360 2508
rect 4068 2456 4120 2508
rect 2872 2388 2924 2440
rect 11612 2524 11664 2576
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 12072 2456 12124 2508
rect 14740 2456 14792 2508
rect 17408 2456 17460 2508
rect 20168 2456 20220 2508
rect 22744 2456 22796 2508
rect 27344 2456 27396 2508
rect 8300 2388 8352 2440
rect 9772 2388 9824 2440
rect 12440 2388 12492 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 22008 2388 22060 2440
rect 25412 2388 25464 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 30748 2388 30800 2440
rect 33416 2388 33468 2440
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 4896 2320 4948 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 2044 24336 2096 24342
rect 2044 24278 2096 24284
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1412 19961 1440 21422
rect 1780 20466 1808 23462
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1872 22642 1900 23258
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1964 22234 1992 23054
rect 1952 22228 2004 22234
rect 1952 22170 2004 22176
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1398 19952 1454 19961
rect 1398 19887 1454 19896
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17921 1440 18770
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1872 17814 1900 20878
rect 2056 18306 2084 24278
rect 2240 22778 2268 26200
rect 2778 24440 2834 24449
rect 2778 24375 2834 24384
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2136 21412 2188 21418
rect 2136 21354 2188 21360
rect 1964 18278 2084 18306
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1216 17604 1268 17610
rect 1216 17546 1268 17552
rect 1228 17105 1256 17546
rect 1766 17368 1822 17377
rect 1766 17303 1822 17312
rect 1780 17202 1808 17303
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1306 13424 1362 13433
rect 1306 13359 1362 13368
rect 1320 12850 1348 13359
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1308 12232 1360 12238
rect 1306 12200 1308 12209
rect 1360 12200 1362 12209
rect 1306 12135 1362 12144
rect 1320 11898 1348 12135
rect 1308 11892 1360 11898
rect 1308 11834 1360 11840
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 6497 1348 6666
rect 1412 6662 1440 15263
rect 1766 13968 1822 13977
rect 1766 13903 1768 13912
rect 1820 13903 1822 13912
rect 1768 13874 1820 13880
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12782 1900 13126
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1674 12608 1730 12617
rect 1674 12543 1730 12552
rect 1688 12434 1716 12543
rect 1688 12406 1900 12434
rect 1582 11792 1638 11801
rect 1582 11727 1638 11736
rect 1596 10130 1624 11727
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1596 10010 1624 10066
rect 1504 9982 1624 10010
rect 1504 9722 1532 9982
rect 1582 9752 1638 9761
rect 1492 9716 1544 9722
rect 1582 9687 1638 9696
rect 1492 9658 1544 9664
rect 1596 9654 1624 9687
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1596 9042 1624 9590
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1688 8090 1716 9454
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1780 6798 1808 8871
rect 1872 7410 1900 12406
rect 1964 12170 1992 18278
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2056 17513 2084 18158
rect 2042 17504 2098 17513
rect 2042 17439 2098 17448
rect 2042 16144 2098 16153
rect 2042 16079 2098 16088
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 7546 1992 11630
rect 2056 7546 2084 16079
rect 2148 11694 2176 21354
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2240 9586 2268 21490
rect 2332 11762 2360 24142
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2412 22500 2464 22506
rect 2412 22442 2464 22448
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2424 10674 2452 22442
rect 2608 14113 2636 23666
rect 2792 23526 2820 24375
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2884 23186 2912 26200
rect 3330 25664 3386 25673
rect 3330 25599 3386 25608
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22250 2820 22986
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3252 22001 3280 22034
rect 3238 21992 3294 22001
rect 3238 21927 3294 21936
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2792 19530 2820 20334
rect 2884 19938 2912 20810
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2884 19910 3004 19938
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2700 19502 2820 19530
rect 2700 19145 2728 19502
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2686 19136 2742 19145
rect 2686 19071 2742 19080
rect 2792 18329 2820 19314
rect 2884 18737 2912 19722
rect 2976 19553 3004 19910
rect 2962 19544 3018 19553
rect 2962 19479 3018 19488
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2870 18728 2926 18737
rect 2870 18663 2926 18672
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2686 18184 2742 18193
rect 2686 18119 2742 18128
rect 2594 14104 2650 14113
rect 2594 14039 2650 14048
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2516 12434 2544 13806
rect 2516 12406 2636 12434
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2516 11218 2544 12106
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2608 9518 2636 12406
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2502 9344 2558 9353
rect 2502 9279 2558 9288
rect 2410 8120 2466 8129
rect 2410 8055 2466 8064
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 2424 6798 2452 8055
rect 2516 7410 2544 9279
rect 2700 9178 2728 18119
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2870 16688 2926 16697
rect 2870 16623 2926 16632
rect 2778 13832 2834 13841
rect 2778 13767 2834 13776
rect 2792 13394 2820 13767
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2884 12442 2912 16623
rect 3344 16182 3372 25599
rect 3528 24274 3556 26200
rect 4066 25256 4122 25265
rect 4066 25191 4122 25200
rect 4080 24954 4108 25191
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 3606 24848 3662 24857
rect 3606 24783 3662 24792
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3620 24070 3648 24783
rect 3608 24064 3660 24070
rect 3514 24032 3570 24041
rect 3608 24006 3660 24012
rect 3514 23967 3570 23976
rect 3528 23866 3556 23967
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 4172 23798 4200 26200
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3700 22976 3752 22982
rect 3700 22918 3752 22924
rect 3712 22710 3740 22918
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 21894 3464 22510
rect 3514 22128 3570 22137
rect 3514 22063 3570 22072
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3436 21146 3464 21830
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3436 15994 3464 21082
rect 3528 19446 3556 22063
rect 3620 20641 3648 22578
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3606 20632 3662 20641
rect 3606 20567 3662 20576
rect 3606 20496 3662 20505
rect 3606 20431 3662 20440
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3620 19258 3648 20431
rect 3712 19718 3740 22374
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3528 19230 3648 19258
rect 3528 17762 3556 19230
rect 3606 17912 3662 17921
rect 3606 17847 3608 17856
rect 3660 17847 3662 17856
rect 3608 17818 3660 17824
rect 3528 17734 3648 17762
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3344 15966 3464 15994
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 3344 13954 3372 15966
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3436 14074 3464 15438
rect 3528 15162 3556 16050
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3514 14920 3570 14929
rect 3620 14890 3648 17734
rect 3514 14855 3570 14864
rect 3608 14884 3660 14890
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3344 13926 3464 13954
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3330 13288 3386 13297
rect 3330 13223 3332 13232
rect 3384 13223 3386 13232
rect 3332 13194 3384 13200
rect 3436 12782 3464 13926
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 11286 2820 11630
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 3330 11248 3386 11257
rect 3330 11183 3386 11192
rect 2778 10976 2834 10985
rect 2778 10911 2834 10920
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2792 8498 2820 10911
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2884 8974 2912 10095
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3344 8634 3372 11183
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 2870 8528 2926 8537
rect 2780 8492 2832 8498
rect 3344 8498 3372 8570
rect 2870 8463 2926 8472
rect 3332 8492 3384 8498
rect 2780 8434 2832 8440
rect 2884 7886 2912 8463
rect 3332 8434 3384 8440
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 3436 8090 3464 11290
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 3436 7818 3464 8026
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3528 7546 3556 14855
rect 3608 14826 3660 14832
rect 3606 13016 3662 13025
rect 3606 12951 3662 12960
rect 3620 11354 3648 12951
rect 3712 12918 3740 19314
rect 3804 17218 3832 23666
rect 4066 23624 4122 23633
rect 4264 23610 4292 24142
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 4066 23559 4068 23568
rect 4120 23559 4122 23568
rect 4172 23582 4292 23610
rect 4068 23530 4120 23536
rect 4066 23216 4122 23225
rect 4066 23151 4122 23160
rect 3976 23044 4028 23050
rect 3976 22986 4028 22992
rect 3882 22808 3938 22817
rect 3882 22743 3938 22752
rect 3896 20534 3924 22743
rect 3988 22506 4016 22986
rect 4080 22710 4108 23151
rect 4172 23118 4200 23582
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 4068 22568 4120 22574
rect 4172 22545 4200 23054
rect 4068 22510 4120 22516
rect 4158 22536 4214 22545
rect 3976 22500 4028 22506
rect 3976 22442 4028 22448
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3988 22030 4016 22102
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3974 21176 4030 21185
rect 3974 21111 4030 21120
rect 3988 21010 4016 21111
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4080 20618 4108 22510
rect 4158 22471 4214 22480
rect 4356 21622 4384 23122
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4344 21616 4396 21622
rect 4344 21558 4396 21564
rect 4250 21040 4306 21049
rect 4250 20975 4252 20984
rect 4304 20975 4306 20984
rect 4252 20946 4304 20952
rect 3988 20590 4108 20618
rect 4344 20596 4396 20602
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3988 18970 4016 20590
rect 4344 20538 4396 20544
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3896 17882 3924 18566
rect 3988 18426 4016 18566
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 4080 18306 4108 20402
rect 4356 20058 4384 20538
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 3988 18278 4108 18306
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3804 17190 3924 17218
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3804 12850 3832 16050
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3606 11248 3662 11257
rect 3606 11183 3608 11192
rect 3660 11183 3662 11192
rect 3608 11154 3660 11160
rect 3620 10810 3648 11154
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3606 10568 3662 10577
rect 3606 10503 3662 10512
rect 3620 9738 3648 10503
rect 3712 10130 3740 12718
rect 3804 10266 3832 12786
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3896 10130 3924 17190
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 3620 9710 3740 9738
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3620 9450 3648 9551
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3712 7954 3740 9710
rect 3804 9586 3832 9930
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3988 8634 4016 18278
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4080 15162 4108 15982
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4066 15056 4122 15065
rect 4172 15026 4200 17614
rect 4066 14991 4068 15000
rect 4120 14991 4122 15000
rect 4160 15020 4212 15026
rect 4068 14962 4120 14968
rect 4160 14962 4212 14968
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4080 11694 4108 14826
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4172 14362 4200 14554
rect 4264 14482 4292 19654
rect 4448 18358 4476 22714
rect 4540 19378 4568 23054
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4540 18766 4568 19178
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4434 17776 4490 17785
rect 4434 17711 4490 17720
rect 4344 17604 4396 17610
rect 4344 17546 4396 17552
rect 4356 16998 4384 17546
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4172 14334 4292 14362
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14074 4200 14214
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4264 14006 4292 14334
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 4250 13560 4306 13569
rect 4250 13495 4306 13504
rect 4158 12472 4214 12481
rect 4158 12407 4214 12416
rect 4172 12238 4200 12407
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4264 11286 4292 13495
rect 4356 12918 4384 15302
rect 4448 15065 4476 17711
rect 4632 17678 4660 18702
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4724 17218 4752 22918
rect 4816 18698 4844 23122
rect 5000 22094 5028 23802
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26330 7434 27000
rect 8022 26330 8078 27000
rect 7116 26302 7434 26330
rect 5460 23662 5488 26200
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5000 22066 5120 22094
rect 4896 21412 4948 21418
rect 4896 21354 4948 21360
rect 4908 19514 4936 21354
rect 5092 20210 5120 22066
rect 5000 20182 5120 20210
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 17882 4844 18634
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4632 17190 4752 17218
rect 4526 16552 4582 16561
rect 4526 16487 4582 16496
rect 4434 15056 4490 15065
rect 4434 14991 4490 15000
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14482 4476 14758
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4448 13258 4476 14418
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4356 12442 4384 12854
rect 4448 12850 4476 13194
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4540 12306 4568 16487
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4068 10056 4120 10062
rect 4066 10024 4068 10033
rect 4120 10024 4122 10033
rect 4066 9959 4122 9968
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4172 8090 4200 8434
rect 4356 8362 4384 12174
rect 4540 11642 4568 12242
rect 4448 11614 4568 11642
rect 4448 10062 4476 11614
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4526 9616 4582 9625
rect 4526 9551 4582 9560
rect 4540 9518 4568 9551
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4632 9178 4660 17190
rect 4710 16824 4766 16833
rect 4710 16759 4766 16768
rect 4724 15348 4752 16759
rect 4908 16250 4936 19314
rect 5000 17270 5028 20182
rect 5184 20074 5212 23190
rect 5092 20046 5212 20074
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 5092 16402 5120 20046
rect 5276 19938 5304 23462
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 5184 19910 5304 19938
rect 5184 16522 5212 19910
rect 5368 19417 5396 22646
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5552 21434 5580 21626
rect 5828 21622 5856 21830
rect 5816 21616 5868 21622
rect 5630 21584 5686 21593
rect 5816 21558 5868 21564
rect 5630 21519 5632 21528
rect 5684 21519 5686 21528
rect 5632 21490 5684 21496
rect 5552 21406 5764 21434
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5460 20058 5488 20878
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5354 19408 5410 19417
rect 5354 19343 5410 19352
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5368 18222 5396 18906
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5368 17241 5396 18158
rect 5354 17232 5410 17241
rect 5354 17167 5410 17176
rect 5172 16516 5224 16522
rect 5368 16504 5396 17167
rect 5460 16697 5488 19110
rect 5446 16688 5502 16697
rect 5446 16623 5502 16632
rect 5368 16476 5488 16504
rect 5172 16458 5224 16464
rect 5092 16374 5396 16402
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 4804 15360 4856 15366
rect 4724 15320 4804 15348
rect 4804 15302 4856 15308
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4724 14618 4752 15030
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4710 13696 4766 13705
rect 4710 13631 4766 13640
rect 4724 12442 4752 13631
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4816 12238 4844 15302
rect 5184 14657 5212 15302
rect 5170 14648 5226 14657
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4988 14612 5040 14618
rect 5170 14583 5226 14592
rect 4988 14554 5040 14560
rect 4908 13870 4936 14554
rect 5000 14074 5028 14554
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 5000 12986 5028 14010
rect 5184 13530 5212 14350
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5184 13394 5212 13466
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5184 12306 5212 13330
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 5276 11762 5304 13670
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 4986 11520 5042 11529
rect 4986 11455 5042 11464
rect 4894 11384 4950 11393
rect 4894 11319 4950 11328
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3698 7712 3754 7721
rect 3698 7647 3754 7656
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 3344 7342 3372 7482
rect 3712 7410 3740 7647
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 2780 7336 2832 7342
rect 3332 7336 3384 7342
rect 2780 7278 2832 7284
rect 2870 7304 2926 7313
rect 2792 6934 2820 7278
rect 3332 7278 3384 7284
rect 2870 7239 2926 7248
rect 2780 6928 2832 6934
rect 2778 6896 2780 6905
rect 2832 6896 2834 6905
rect 2778 6831 2834 6840
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1306 6488 1362 6497
rect 1780 6458 1808 6734
rect 1306 6423 1362 6432
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 2884 6322 2912 7239
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3988 6458 4016 6598
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1320 6089 1348 6190
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1320 5914 1348 6015
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 1360 5672 1362 5681
rect 1306 5607 1362 5616
rect 1306 5264 1362 5273
rect 1306 5199 1308 5208
rect 1360 5199 1362 5208
rect 1308 5170 1360 5176
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 1306 4856 1362 4865
rect 2950 4859 3258 4868
rect 1306 4791 1362 4800
rect 1320 4690 1348 4791
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 2780 4480 2832 4486
rect 1766 4448 1822 4457
rect 2780 4422 2832 4428
rect 3514 4448 3570 4457
rect 1766 4383 1822 4392
rect 1780 4146 1808 4383
rect 2792 4214 2820 4422
rect 3514 4383 3570 4392
rect 2780 4208 2832 4214
rect 2686 4176 2742 4185
rect 1768 4140 1820 4146
rect 2780 4150 2832 4156
rect 2686 4111 2742 4120
rect 1768 4082 1820 4088
rect 2700 4010 2728 4111
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2792 3738 2820 4150
rect 3528 4146 3556 4383
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 2884 4049 2912 4082
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 1308 3732 1360 3738
rect 1308 3674 1360 3680
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 1320 3641 1348 3674
rect 1306 3632 1362 3641
rect 1306 3567 1362 3576
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3233 1348 3470
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1320 2825 1348 2926
rect 1400 2848 1452 2854
rect 1306 2816 1362 2825
rect 1400 2790 1452 2796
rect 1306 2751 1362 2760
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1320 2417 1348 2450
rect 1306 2408 1362 2417
rect 1306 2343 1362 2352
rect 1412 800 1440 2790
rect 2792 2009 2820 2994
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2446 2912 2790
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 3344 1601 3372 3334
rect 3436 3194 3464 3402
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 4080 800 4108 2450
rect 4908 2378 4936 11319
rect 5000 10606 5028 11455
rect 5368 10674 5396 16374
rect 5460 13870 5488 16476
rect 5552 15570 5580 21286
rect 5630 19952 5686 19961
rect 5630 19887 5686 19896
rect 5644 18290 5672 19887
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 17921 5672 18226
rect 5630 17912 5686 17921
rect 5630 17847 5686 17856
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5644 15910 5672 17138
rect 5736 16794 5764 21406
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5828 17134 5856 20334
rect 5920 17252 5948 23530
rect 6012 18222 6040 24006
rect 6104 23186 6132 26200
rect 6644 24200 6696 24206
rect 6550 24168 6606 24177
rect 6748 24188 6776 26200
rect 7012 25560 7064 25566
rect 7012 25502 7064 25508
rect 6748 24160 6868 24188
rect 6644 24142 6696 24148
rect 6550 24103 6606 24112
rect 6564 24070 6592 24103
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6104 20466 6132 21830
rect 6196 21593 6224 23462
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6182 21584 6238 21593
rect 6182 21519 6238 21528
rect 6288 20777 6316 23054
rect 6656 22642 6684 24142
rect 6736 23520 6788 23526
rect 6734 23488 6736 23497
rect 6788 23488 6790 23497
rect 6734 23423 6790 23432
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6380 21350 6408 22374
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6380 20806 6408 21286
rect 6368 20800 6420 20806
rect 6274 20768 6330 20777
rect 6368 20742 6420 20748
rect 6274 20703 6330 20712
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5920 17224 6040 17252
rect 5816 17128 5868 17134
rect 5908 17128 5960 17134
rect 5816 17070 5868 17076
rect 5906 17096 5908 17105
rect 5960 17096 5962 17105
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5828 16182 5856 17070
rect 5906 17031 5962 17040
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5632 15904 5684 15910
rect 5736 15881 5764 15982
rect 5632 15846 5684 15852
rect 5722 15872 5778 15881
rect 5722 15807 5778 15816
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5538 14784 5594 14793
rect 5538 14719 5594 14728
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 9586 5212 10406
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5276 8634 5304 10610
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5368 8566 5396 10503
rect 5460 9674 5488 13670
rect 5552 12170 5580 14719
rect 5722 14512 5778 14521
rect 5722 14447 5778 14456
rect 5632 13932 5684 13938
rect 5736 13920 5764 14447
rect 5828 14346 5856 14962
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5920 14226 5948 17031
rect 5684 13892 5764 13920
rect 5632 13874 5684 13880
rect 5736 12986 5764 13892
rect 5828 14198 5948 14226
rect 5828 13734 5856 14198
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5920 13190 5948 13738
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5644 11898 5672 12582
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5632 11688 5684 11694
rect 5736 11642 5764 12106
rect 5684 11636 5764 11642
rect 5632 11630 5764 11636
rect 5540 11620 5592 11626
rect 5644 11614 5764 11630
rect 5540 11562 5592 11568
rect 5552 11354 5580 11562
rect 5736 11354 5764 11614
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5828 10130 5856 12854
rect 5920 11694 5948 13126
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5460 9646 5580 9674
rect 6012 9654 6040 17224
rect 6104 16561 6132 20266
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 6196 18630 6224 19722
rect 6380 18630 6408 19858
rect 6472 19514 6500 22374
rect 6656 22137 6684 22578
rect 6642 22128 6698 22137
rect 6642 22063 6698 22072
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 19961 6592 21966
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6550 19952 6606 19961
rect 6550 19887 6606 19896
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6458 19408 6514 19417
rect 6458 19343 6460 19352
rect 6512 19343 6514 19352
rect 6552 19372 6604 19378
rect 6460 19314 6512 19320
rect 6552 19314 6604 19320
rect 6564 19174 6592 19314
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6196 17610 6224 18566
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6288 17921 6316 18226
rect 6274 17912 6330 17921
rect 6274 17847 6330 17856
rect 6184 17604 6236 17610
rect 6184 17546 6236 17552
rect 6196 17202 6224 17546
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16794 6224 16934
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6090 16552 6146 16561
rect 6090 16487 6146 16496
rect 6288 16436 6316 17847
rect 6550 17640 6606 17649
rect 6550 17575 6606 17584
rect 6458 17368 6514 17377
rect 6458 17303 6514 17312
rect 6472 17270 6500 17303
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6104 16408 6316 16436
rect 5552 8974 5580 9646
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5172 8560 5224 8566
rect 5000 8508 5172 8514
rect 5000 8502 5224 8508
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5000 8498 5212 8502
rect 4988 8492 5212 8498
rect 5040 8486 5212 8492
rect 4988 8434 5040 8440
rect 6104 7750 6132 16408
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6196 15638 6224 15982
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6196 15065 6224 15574
rect 6380 15450 6408 17138
rect 6564 17105 6592 17575
rect 6550 17096 6606 17105
rect 6550 17031 6606 17040
rect 6458 16688 6514 16697
rect 6458 16623 6514 16632
rect 6288 15422 6408 15450
rect 6288 15094 6316 15422
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6276 15088 6328 15094
rect 6182 15056 6238 15065
rect 6276 15030 6328 15036
rect 6182 14991 6184 15000
rect 6236 14991 6238 15000
rect 6184 14962 6236 14968
rect 6288 14346 6316 15030
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6288 13938 6316 14282
rect 6380 14074 6408 15302
rect 6472 15178 6500 16623
rect 6656 16130 6684 21422
rect 6748 17066 6776 22578
rect 6840 21962 6868 24160
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6932 23526 6960 23598
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6840 18170 6868 20334
rect 6932 19446 6960 22714
rect 7024 21350 7052 25502
rect 7116 24274 7144 26302
rect 7378 26200 7434 26302
rect 7852 26302 8078 26330
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 7208 23633 7236 24142
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7194 23624 7250 23633
rect 7194 23559 7250 23568
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 22166 7144 22374
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 7024 20942 7052 21286
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7116 20754 7144 21966
rect 7024 20726 7144 20754
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6918 19272 6974 19281
rect 6918 19207 6974 19216
rect 6932 18290 6960 19207
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6840 18142 6960 18170
rect 6932 18086 6960 18142
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6748 16561 6776 16594
rect 6734 16552 6790 16561
rect 6734 16487 6790 16496
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6564 16102 6684 16130
rect 6564 16046 6592 16102
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6550 15872 6606 15881
rect 6550 15807 6606 15816
rect 6564 15348 6592 15807
rect 6656 15609 6684 15982
rect 6642 15600 6698 15609
rect 6642 15535 6698 15544
rect 6564 15320 6684 15348
rect 6472 15150 6592 15178
rect 6564 14362 6592 15150
rect 6472 14334 6592 14362
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6288 13530 6316 13874
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6288 13326 6316 13466
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6288 13190 6316 13262
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12170 6316 13126
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6288 11132 6316 12106
rect 6368 11144 6420 11150
rect 6182 11112 6238 11121
rect 6288 11104 6368 11132
rect 6368 11086 6420 11092
rect 6182 11047 6238 11056
rect 6196 9042 6224 11047
rect 6366 10432 6422 10441
rect 6366 10367 6422 10376
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6380 8498 6408 10367
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6472 8430 6500 14334
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6564 11762 6592 12922
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6656 8838 6684 15320
rect 6748 14482 6776 16390
rect 6840 15570 6868 18022
rect 6932 16454 6960 18022
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6932 15450 6960 15506
rect 6840 15422 6960 15450
rect 6840 14822 6868 15422
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6932 13258 6960 15098
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 7024 12918 7052 20726
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7116 17678 7144 20198
rect 7208 19310 7236 20742
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7208 18358 7236 19246
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7194 18048 7250 18057
rect 7194 17983 7250 17992
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7208 17490 7236 17983
rect 7116 17462 7236 17490
rect 7116 12986 7144 17462
rect 7300 17320 7328 23734
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 21146 7420 22510
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7392 21010 7420 21082
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7484 20754 7512 24890
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7576 21622 7604 23598
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7392 20466 7420 20742
rect 7484 20726 7604 20754
rect 7380 20460 7432 20466
rect 7432 20420 7512 20448
rect 7380 20402 7432 20408
rect 7380 20324 7432 20330
rect 7380 20266 7432 20272
rect 7392 18154 7420 20266
rect 7484 19786 7512 20420
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7576 19446 7604 20726
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7576 17610 7604 18906
rect 7668 17882 7696 22578
rect 7760 21894 7788 23462
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 21616 7892 21622
rect 7840 21558 7892 21564
rect 7852 19718 7880 21558
rect 8312 21350 8340 23054
rect 8484 23044 8536 23050
rect 8484 22986 8536 22992
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8114 20904 8170 20913
rect 8114 20839 8170 20848
rect 8128 20806 8156 20839
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20058 8340 21286
rect 8404 20874 8432 21830
rect 8496 21010 8524 22986
rect 8680 22574 8708 26200
rect 9126 24848 9182 24857
rect 9126 24783 9182 24792
rect 9140 24070 9168 24783
rect 9324 24342 9352 26200
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9876 23730 9904 25094
rect 9968 23798 9996 26200
rect 10140 25628 10192 25634
rect 10140 25570 10192 25576
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10060 24206 10088 25298
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8666 21584 8722 21593
rect 8666 21519 8722 21528
rect 8680 21146 8708 21519
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7760 19094 8156 19122
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 7380 17332 7432 17338
rect 7300 17292 7380 17320
rect 7380 17274 7432 17280
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7208 15706 7236 17138
rect 7484 16998 7512 17546
rect 7576 17134 7604 17546
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7484 16561 7512 16934
rect 7576 16794 7604 16934
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7656 16584 7708 16590
rect 7470 16552 7526 16561
rect 7656 16526 7708 16532
rect 7470 16487 7526 16496
rect 7668 16402 7696 16526
rect 7760 16522 7788 19094
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7852 17746 7880 18906
rect 8128 18902 8156 19094
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7944 17592 7972 17750
rect 7852 17564 7972 17592
rect 7852 16998 7880 17564
rect 8312 17542 8340 19654
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8496 18204 8524 18770
rect 8588 18630 8616 21082
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8576 18216 8628 18222
rect 8496 18176 8576 18204
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7668 16374 7788 16402
rect 7380 16244 7432 16250
rect 7300 16204 7380 16232
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7196 15496 7248 15502
rect 7194 15464 7196 15473
rect 7248 15464 7250 15473
rect 7194 15399 7250 15408
rect 7208 14550 7236 15399
rect 7300 14958 7328 16204
rect 7380 16186 7432 16192
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7102 12880 7158 12889
rect 6920 12844 6972 12850
rect 7102 12815 7158 12824
rect 6920 12786 6972 12792
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 11830 6868 12582
rect 6932 12434 6960 12786
rect 6932 12406 7052 12434
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 11014 6776 11086
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10742 6776 10950
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6748 10266 6776 10678
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6840 10130 6868 11154
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9110 6868 9454
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6932 8362 6960 12038
rect 7024 11626 7052 12406
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 7010 11520 7066 11529
rect 7010 11455 7066 11464
rect 7024 10674 7052 11455
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 8514 7052 10474
rect 7116 9586 7144 12815
rect 7208 12617 7236 14350
rect 7300 14074 7328 14758
rect 7392 14074 7420 16050
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7484 15366 7512 15982
rect 7562 15736 7618 15745
rect 7562 15671 7618 15680
rect 7576 15638 7604 15671
rect 7564 15632 7616 15638
rect 7564 15574 7616 15580
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13258 7328 13806
rect 7484 13734 7512 15302
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7194 12608 7250 12617
rect 7194 12543 7250 12552
rect 7300 12374 7328 13194
rect 7392 12646 7420 13330
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7392 11762 7420 12582
rect 7576 12434 7604 15370
rect 7668 15337 7696 16050
rect 7654 15328 7710 15337
rect 7654 15263 7710 15272
rect 7760 15094 7788 16374
rect 7852 15366 7880 16934
rect 8022 16824 8078 16833
rect 8022 16759 8024 16768
rect 8076 16759 8078 16768
rect 8024 16730 8076 16736
rect 8128 16697 8156 17274
rect 8114 16688 8170 16697
rect 8114 16623 8170 16632
rect 8128 16590 8156 16623
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16232 8340 17478
rect 8404 17338 8432 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8220 16204 8340 16232
rect 8220 16046 8248 16204
rect 8404 16153 8432 17138
rect 8390 16144 8446 16153
rect 8300 16108 8352 16114
rect 8496 16114 8524 18176
rect 8576 18158 8628 18164
rect 8390 16079 8446 16088
rect 8484 16108 8536 16114
rect 8300 16050 8352 16056
rect 8484 16050 8536 16056
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8312 15570 8340 16050
rect 8482 16008 8538 16017
rect 8482 15943 8538 15952
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7838 15056 7894 15065
rect 7656 14952 7708 14958
rect 7654 14920 7656 14929
rect 7708 14920 7710 14929
rect 7654 14855 7710 14864
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7668 13938 7696 14486
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 13190 7696 13738
rect 7760 13530 7788 15030
rect 7838 14991 7894 15000
rect 7852 14958 7880 14991
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 14414 7880 14894
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7484 12406 7604 12434
rect 7484 12238 7512 12406
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 9994 7236 11630
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7286 10704 7342 10713
rect 7286 10639 7342 10648
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7208 9382 7236 9930
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7194 9208 7250 9217
rect 7194 9143 7196 9152
rect 7248 9143 7250 9152
rect 7196 9114 7248 9120
rect 7300 8634 7328 10639
rect 7392 10606 7420 11562
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 9722 7420 10406
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7392 8514 7420 8570
rect 7024 8486 7420 8514
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6274 4176 6330 4185
rect 6274 4111 6276 4120
rect 6328 4111 6330 4120
rect 6276 4082 6328 4088
rect 6932 3126 6960 8298
rect 7024 3602 7052 8486
rect 7484 6186 7512 12174
rect 7668 11830 7696 13126
rect 7760 12714 7788 13330
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7746 12608 7802 12617
rect 7746 12543 7802 12552
rect 7760 12306 7788 12543
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7852 11642 7880 14214
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8220 12238 8248 12310
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8208 11824 8260 11830
rect 8206 11792 8208 11801
rect 8260 11792 8262 11801
rect 8206 11727 8262 11736
rect 8116 11688 8168 11694
rect 7852 11614 7972 11642
rect 8116 11630 8168 11636
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7576 9994 7604 10202
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7668 7342 7696 11494
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7760 9518 7788 11222
rect 7852 10470 7880 11494
rect 7944 11082 7972 11614
rect 8128 11218 8156 11630
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 8220 11014 8248 11727
rect 8312 11150 8340 14826
rect 8496 12434 8524 15943
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8588 15094 8616 15846
rect 8680 15706 8708 19314
rect 8772 18834 8800 23666
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 22778 9076 22918
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 9220 22092 9272 22098
rect 9220 22034 9272 22040
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8772 17134 8800 18634
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 16454 8800 16934
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8666 15600 8722 15609
rect 8666 15535 8722 15544
rect 8680 15502 8708 15535
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8680 15162 8708 15302
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8772 14793 8800 16390
rect 8864 15094 8892 22034
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21622 8984 21830
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8956 20466 8984 21558
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 9048 19922 9076 20198
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 17202 9076 18770
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9140 17610 9168 18090
rect 9232 18057 9260 22034
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9218 18048 9274 18057
rect 9218 17983 9274 17992
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 9034 17096 9090 17105
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 8956 14906 8984 17070
rect 9034 17031 9090 17040
rect 9048 16998 9076 17031
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9048 15094 9076 16458
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 8864 14878 8984 14906
rect 8758 14784 8814 14793
rect 8758 14719 8814 14728
rect 8574 14648 8630 14657
rect 8574 14583 8630 14592
rect 8588 14006 8616 14583
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8404 12406 8524 12434
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8208 11008 8260 11014
rect 8260 10968 8340 10996
rect 8208 10950 8260 10956
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8312 10742 8340 10968
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 10130 7880 10406
rect 8128 10198 8156 10542
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 9586 7880 10066
rect 8220 10010 8248 10406
rect 8220 9982 8340 10010
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8312 9602 8340 9982
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7944 9574 8340 9602
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7746 9072 7802 9081
rect 7746 9007 7802 9016
rect 7760 8974 7788 9007
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8498 7788 8910
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7852 3058 7880 9522
rect 7944 8974 7972 9574
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8312 8090 8340 8774
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 8022 8432 12406
rect 8588 8498 8616 12854
rect 8680 10554 8708 14418
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13258 8800 14214
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 12918 8800 13194
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8772 11801 8800 12854
rect 8758 11792 8814 11801
rect 8758 11727 8814 11736
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 11286 8800 11494
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8760 10600 8812 10606
rect 8680 10548 8760 10554
rect 8680 10542 8812 10548
rect 8680 10526 8800 10542
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8680 9110 8708 9590
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8772 9042 8800 9318
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8864 6866 8892 14878
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8956 12102 8984 13670
rect 9048 13394 9076 13670
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 9048 11626 9076 12718
rect 9140 12170 9168 17546
rect 9218 15600 9274 15609
rect 9218 15535 9220 15544
rect 9272 15535 9274 15544
rect 9220 15506 9272 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 14618 9260 15370
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9048 11286 9076 11562
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9232 11218 9260 14010
rect 9324 13954 9352 20878
rect 9416 20505 9444 21830
rect 9508 21690 9536 21966
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9600 21622 9628 22986
rect 10152 22642 10180 25570
rect 10704 22710 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10784 25084 10836 25090
rect 10784 25026 10836 25032
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10796 22556 10824 25026
rect 10704 22528 10824 22556
rect 9784 22222 10088 22250
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9692 21894 9720 22102
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9784 21690 9812 22222
rect 10060 22030 10088 22222
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9784 21350 9812 21490
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9772 21344 9824 21350
rect 9770 21312 9772 21321
rect 9824 21312 9826 21321
rect 9770 21247 9826 21256
rect 9402 20496 9458 20505
rect 9402 20431 9458 20440
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9416 20058 9444 20334
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9416 17746 9444 19994
rect 9692 19310 9720 20334
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9876 18986 9904 21422
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9968 19446 9996 20470
rect 10152 20262 10180 22034
rect 10230 21448 10286 21457
rect 10230 21383 10232 21392
rect 10284 21383 10286 21392
rect 10232 21354 10284 21360
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10612 20806 10640 21014
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9692 18958 9904 18986
rect 9494 18456 9550 18465
rect 9494 18391 9550 18400
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9508 17082 9536 18391
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 17921 9628 18158
rect 9586 17912 9642 17921
rect 9586 17847 9642 17856
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9416 17054 9536 17082
rect 9416 14346 9444 17054
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 15745 9536 16934
rect 9494 15736 9550 15745
rect 9494 15671 9550 15680
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9508 14521 9536 14826
rect 9494 14512 9550 14521
rect 9494 14447 9550 14456
rect 9600 14362 9628 17138
rect 9692 15881 9720 18958
rect 9770 18864 9826 18873
rect 9770 18799 9826 18808
rect 10048 18828 10100 18834
rect 9784 18358 9812 18799
rect 10048 18770 10100 18776
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9784 17338 9812 18294
rect 9968 17746 9996 18634
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9954 17368 10010 17377
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9864 17332 9916 17338
rect 9954 17303 10010 17312
rect 9864 17274 9916 17280
rect 9770 17232 9826 17241
rect 9876 17202 9904 17274
rect 9968 17202 9996 17303
rect 9770 17167 9826 17176
rect 9864 17196 9916 17202
rect 9784 17066 9812 17167
rect 9864 17138 9916 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9678 15872 9734 15881
rect 9678 15807 9734 15816
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9508 14334 9628 14362
rect 9692 14346 9720 14418
rect 9784 14414 9812 16390
rect 9876 16017 9904 17138
rect 10060 16232 10088 18770
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10152 16590 10180 18702
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10244 18086 10272 18634
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10336 17882 10364 19450
rect 10428 19417 10456 19450
rect 10414 19408 10470 19417
rect 10414 19343 10470 19352
rect 10520 18902 10548 19790
rect 10704 19446 10732 22528
rect 10888 22488 10916 25434
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 10796 22460 10916 22488
rect 10796 22030 10824 22460
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 11164 21554 11192 22986
rect 11256 22098 11284 26200
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11716 24410 11744 24754
rect 11900 24426 11928 26200
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 11704 24404 11756 24410
rect 11900 24398 12020 24426
rect 11704 24346 11756 24352
rect 11886 24304 11942 24313
rect 11886 24239 11942 24248
rect 11900 24206 11928 24239
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11520 23520 11572 23526
rect 11888 23520 11940 23526
rect 11520 23462 11572 23468
rect 11886 23488 11888 23497
rect 11940 23488 11942 23497
rect 11532 23050 11560 23462
rect 11886 23423 11942 23432
rect 11520 23044 11572 23050
rect 11888 23044 11940 23050
rect 11572 23004 11888 23032
rect 11520 22986 11572 22992
rect 11888 22986 11940 22992
rect 11794 22808 11850 22817
rect 11794 22743 11850 22752
rect 11808 22710 11836 22743
rect 11900 22710 11928 22986
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11440 21950 11652 21978
rect 11808 21962 11836 22646
rect 11992 22166 12020 24398
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11440 21894 11468 21950
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11164 20942 11192 21490
rect 11242 21448 11298 21457
rect 11242 21383 11298 21392
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11164 20534 11192 20878
rect 11152 20528 11204 20534
rect 11072 20488 11152 20516
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10888 20058 10916 20198
rect 11072 20058 11100 20488
rect 11152 20470 11204 20476
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11072 19854 11100 19994
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10980 19514 11008 19722
rect 11164 19718 11192 20334
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10692 19440 10744 19446
rect 10744 19388 10824 19394
rect 10692 19382 10824 19388
rect 10704 19366 10824 19382
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16250 10180 16526
rect 10244 16250 10272 17614
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 9968 16204 10088 16232
rect 10140 16244 10192 16250
rect 9968 16046 9996 16204
rect 10140 16186 10192 16192
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10046 16144 10102 16153
rect 10046 16079 10102 16088
rect 9956 16040 10008 16046
rect 9862 16008 9918 16017
rect 9956 15982 10008 15988
rect 9862 15943 9918 15952
rect 9862 15464 9918 15473
rect 9862 15399 9864 15408
rect 9916 15399 9918 15408
rect 9956 15428 10008 15434
rect 9864 15370 9916 15376
rect 9956 15370 10008 15376
rect 9862 15192 9918 15201
rect 9862 15127 9918 15136
rect 9876 15094 9904 15127
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9968 15026 9996 15370
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 14550 9904 14894
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14340 9732 14346
rect 9324 13926 9444 13954
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 12646 9352 13806
rect 9416 13734 9444 13926
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9508 13569 9536 14334
rect 9680 14282 9732 14288
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9494 13560 9550 13569
rect 9494 13495 9550 13504
rect 9402 13424 9458 13433
rect 9402 13359 9404 13368
rect 9456 13359 9458 13368
rect 9404 13330 9456 13336
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12306 9352 12582
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9508 11150 9536 13126
rect 9600 12918 9628 13194
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9692 12442 9720 13194
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9784 11665 9812 14214
rect 9876 12986 9904 14214
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9968 12866 9996 14962
rect 10060 14906 10088 16079
rect 10060 14878 10180 14906
rect 10048 14816 10100 14822
rect 10046 14784 10048 14793
rect 10100 14784 10102 14793
rect 10046 14719 10102 14728
rect 10152 14550 10180 14878
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10060 13870 10088 14486
rect 10152 14346 10180 14486
rect 10244 14482 10272 16186
rect 10336 16153 10364 17002
rect 10428 16726 10456 18566
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 10428 16454 10456 16662
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10322 16144 10378 16153
rect 10322 16079 10378 16088
rect 10428 16046 10456 16390
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9876 12838 9996 12866
rect 9770 11656 9826 11665
rect 9770 11591 9826 11600
rect 9784 11393 9812 11591
rect 9770 11384 9826 11393
rect 9770 11319 9826 11328
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9496 11144 9548 11150
rect 9310 11112 9366 11121
rect 9496 11086 9548 11092
rect 9310 11047 9366 11056
rect 9404 11076 9456 11082
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10266 9076 10406
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9058 9168 9862
rect 9048 9030 9168 9058
rect 9048 7206 9076 9030
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 7546 9168 8842
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9232 7478 9260 10950
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9324 7410 9352 11047
rect 9404 11018 9456 11024
rect 9416 9042 9444 11018
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 9586 9536 10406
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9508 8906 9536 9522
rect 9692 9178 9720 9522
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9600 8634 9628 8978
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9586 8392 9642 8401
rect 9586 8327 9588 8336
rect 9640 8327 9642 8336
rect 9588 8298 9640 8304
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 9692 3942 9720 8774
rect 9784 5710 9812 11154
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9876 5166 9904 12838
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9968 11762 9996 12106
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9968 10810 9996 11698
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10060 10606 10088 13806
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10152 12986 10180 13466
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10060 9110 10088 10542
rect 10152 9178 10180 12718
rect 10244 11218 10272 14282
rect 10336 12850 10364 15914
rect 10428 15366 10456 15982
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10428 12238 10456 14758
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10520 11558 10548 18226
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 10612 14006 10640 16118
rect 10704 14618 10732 17478
rect 10796 15094 10824 19366
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10966 18728 11022 18737
rect 10966 18663 11022 18672
rect 10874 18592 10930 18601
rect 10874 18527 10930 18536
rect 10888 17678 10916 18527
rect 10980 17678 11008 18663
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11072 17241 11100 19246
rect 11256 18714 11284 21383
rect 11532 21146 11560 21830
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11348 20777 11376 20810
rect 11428 20800 11480 20806
rect 11334 20768 11390 20777
rect 11428 20742 11480 20748
rect 11334 20703 11390 20712
rect 11440 20602 11468 20742
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11256 18686 11468 18714
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11058 17232 11114 17241
rect 10876 17196 10928 17202
rect 11058 17167 11114 17176
rect 11152 17196 11204 17202
rect 10876 17138 10928 17144
rect 11152 17138 11204 17144
rect 10888 16153 10916 17138
rect 11164 16969 11192 17138
rect 11150 16960 11206 16969
rect 11150 16895 11206 16904
rect 11348 16658 11376 18566
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11058 16552 11114 16561
rect 11058 16487 11114 16496
rect 10874 16144 10930 16153
rect 10874 16079 10930 16088
rect 10966 16008 11022 16017
rect 10876 15972 10928 15978
rect 10966 15943 10968 15952
rect 10876 15914 10928 15920
rect 11020 15943 11022 15952
rect 10968 15914 11020 15920
rect 10888 15570 10916 15914
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10980 15434 11008 15642
rect 11072 15434 11100 16487
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 11058 15328 11114 15337
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10796 14618 10824 15030
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10888 14414 10916 15302
rect 11058 15263 11114 15272
rect 10966 15192 11022 15201
rect 10966 15127 11022 15136
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10600 14000 10652 14006
rect 10652 13960 10732 13988
rect 10600 13942 10652 13948
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 13462 10640 13738
rect 10704 13530 10732 13960
rect 10782 13832 10838 13841
rect 10782 13767 10838 13776
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10704 12986 10732 13466
rect 10796 13190 10824 13767
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10690 12880 10746 12889
rect 10690 12815 10692 12824
rect 10744 12815 10746 12824
rect 10692 12786 10744 12792
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10612 11830 10640 12038
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10324 11008 10376 11014
rect 10230 10976 10286 10985
rect 10324 10950 10376 10956
rect 10230 10911 10286 10920
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 9104 10100 9110
rect 10100 9052 10180 9058
rect 10048 9046 10180 9052
rect 10060 9030 10180 9046
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9968 7750 9996 8026
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9968 4010 9996 7686
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7208 2650 7236 2926
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 6748 800 6776 2450
rect 8312 2446 8340 3130
rect 10060 3126 10088 8842
rect 10152 7954 10180 9030
rect 10244 8974 10272 10911
rect 10336 8974 10364 10950
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 10130 10548 10406
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10520 6866 10548 8434
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10612 4146 10640 8366
rect 10704 6730 10732 12038
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10266 10824 10950
rect 10980 10810 11008 15127
rect 11072 14414 11100 15263
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11072 13462 11100 14350
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11164 12986 11192 16050
rect 11256 15162 11284 16390
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11348 15042 11376 16594
rect 11256 15014 11376 15042
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12434 11284 15014
rect 11336 14952 11388 14958
rect 11334 14920 11336 14929
rect 11388 14920 11390 14929
rect 11334 14855 11390 14864
rect 11440 14074 11468 18686
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11532 13954 11560 21082
rect 11624 18970 11652 21950
rect 11796 21956 11848 21962
rect 11716 21916 11796 21944
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11624 17882 11652 18090
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11716 16454 11744 21916
rect 11796 21898 11848 21904
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 21078 11836 21286
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 20058 11836 20402
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11794 19816 11850 19825
rect 11794 19751 11850 19760
rect 11808 19718 11836 19751
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11808 18154 11836 18702
rect 11900 18465 11928 20198
rect 11992 19530 12020 21490
rect 12084 20942 12112 25230
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 12360 23866 12388 24618
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12544 23798 12572 26200
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12636 24206 12664 25162
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12268 23633 12296 23666
rect 12254 23624 12310 23633
rect 12254 23559 12310 23568
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22574 12480 23122
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12176 19854 12204 21626
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12268 21078 12296 21422
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 11992 19502 12112 19530
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11886 18456 11942 18465
rect 11886 18391 11942 18400
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11808 15960 11836 17002
rect 11716 15932 11836 15960
rect 11716 15026 11744 15932
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11164 12406 11284 12434
rect 11348 13926 11560 13954
rect 11058 11248 11114 11257
rect 11058 11183 11114 11192
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10888 9518 10916 10134
rect 10980 9994 11008 10202
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 11072 8362 11100 11183
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11164 7954 11192 12406
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11256 12102 11284 12242
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10062 11284 10542
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9518 11284 9998
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11348 7954 11376 13926
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11532 12434 11560 13806
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11624 12646 11652 12951
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11440 12406 11560 12434
rect 11440 7970 11468 12406
rect 11624 12374 11652 12582
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11218 11560 11562
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11532 9994 11560 10746
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11336 7948 11388 7954
rect 11440 7942 11560 7970
rect 11336 7890 11388 7896
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 11440 3738 11468 7822
rect 11532 4690 11560 7942
rect 11624 7478 11652 9318
rect 11716 8022 11744 14010
rect 11808 14006 11836 15302
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11808 13870 11836 13942
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11808 11694 11836 12242
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11900 10010 11928 18226
rect 11992 17678 12020 19382
rect 11980 17672 12032 17678
rect 12084 17649 12112 19502
rect 12268 18834 12296 20334
rect 12360 19922 12388 21558
rect 12452 21554 12480 22510
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12452 20516 12480 21490
rect 12544 21010 12572 22102
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12636 20618 12664 23666
rect 12820 22030 12848 24822
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13188 22710 13216 22986
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22098 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26330 15162 27000
rect 15028 26302 15162 26330
rect 13832 24138 13860 26200
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14292 24410 14320 24686
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14476 24342 14504 26200
rect 14924 25016 14976 25022
rect 14924 24958 14976 24964
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23254 13768 24006
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22574 13492 22918
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 13464 21486 13492 22510
rect 13832 21622 13860 22986
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13832 21010 13860 21558
rect 13924 21185 13952 24142
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14200 21690 14228 22374
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 13910 21176 13966 21185
rect 13910 21111 13966 21120
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 12636 20590 13768 20618
rect 12532 20528 12584 20534
rect 12452 20488 12532 20516
rect 12452 19990 12480 20488
rect 12532 20470 12584 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12544 19836 12572 20334
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12452 19808 12572 19836
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12360 18737 12388 18838
rect 12346 18728 12402 18737
rect 12346 18663 12402 18672
rect 12452 18329 12480 19808
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12636 18442 12664 19722
rect 12728 19718 12756 20198
rect 12820 19990 12848 20402
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13358 20224 13414 20233
rect 12950 20156 13258 20165
rect 13358 20159 13414 20168
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 20058 13400 20159
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12544 18414 12664 18442
rect 12438 18320 12494 18329
rect 12438 18255 12494 18264
rect 12256 18216 12308 18222
rect 12162 18184 12218 18193
rect 12256 18158 12308 18164
rect 12162 18119 12218 18128
rect 12176 18086 12204 18119
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 11980 17614 12032 17620
rect 12070 17640 12126 17649
rect 11992 16114 12020 17614
rect 12268 17610 12296 18158
rect 12070 17575 12126 17584
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12084 16998 12112 17274
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12268 16726 12296 17546
rect 12544 17338 12572 18414
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12256 16720 12308 16726
rect 12452 16697 12480 16934
rect 12256 16662 12308 16668
rect 12438 16688 12494 16697
rect 12438 16623 12494 16632
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12070 16280 12126 16289
rect 12070 16215 12126 16224
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 12084 15910 12112 16215
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12176 15638 12204 16458
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12072 15632 12124 15638
rect 12070 15600 12072 15609
rect 12164 15632 12216 15638
rect 12124 15600 12126 15609
rect 12164 15574 12216 15580
rect 12070 15535 12126 15544
rect 11978 15056 12034 15065
rect 11978 14991 11980 15000
rect 12032 14991 12034 15000
rect 12072 15020 12124 15026
rect 11980 14962 12032 14968
rect 12072 14962 12124 14968
rect 12084 14793 12112 14962
rect 12268 14958 12296 16118
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12070 14784 12126 14793
rect 12070 14719 12126 14728
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13394 12020 14350
rect 12268 14346 12296 14418
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13938 12112 14010
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 12176 12646 12204 13806
rect 12268 13530 12296 14282
rect 12360 13938 12388 16526
rect 12452 16250 12480 16526
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12544 15450 12572 16934
rect 12452 15422 12572 15450
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12360 13734 12388 13874
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 11992 11558 12020 11727
rect 12084 11558 12112 12038
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 10742 12112 11494
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11808 9982 11928 10010
rect 11808 9926 11836 9982
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11888 9920 11940 9926
rect 11992 9874 12020 10066
rect 11940 9868 12020 9874
rect 11888 9862 12020 9868
rect 11900 9846 12020 9862
rect 11992 9654 12020 9846
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11808 8566 11836 8978
rect 11992 8906 12020 9046
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11900 7546 11928 8842
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11992 3534 12020 7958
rect 12176 6254 12204 12582
rect 12268 12306 12296 13194
rect 12452 12918 12480 15422
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12544 12442 12572 15302
rect 12636 15162 12664 18226
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17610 12756 18090
rect 12820 18086 12848 19722
rect 13464 19310 13492 20266
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13268 19236 13320 19242
rect 13320 19196 13400 19224
rect 13268 19178 13320 19184
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13004 18290 13032 18566
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13280 18154 13308 18566
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17882 13400 19196
rect 13556 18834 13584 20470
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13648 20369 13676 20402
rect 13634 20360 13690 20369
rect 13634 20295 13690 20304
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 20097 13676 20198
rect 13634 20088 13690 20097
rect 13634 20023 13690 20032
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13556 17921 13584 18226
rect 13542 17912 13598 17921
rect 13360 17876 13412 17882
rect 13542 17847 13598 17856
rect 13360 17818 13412 17824
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 16182 12756 17546
rect 12898 17368 12954 17377
rect 12898 17303 12954 17312
rect 12912 17270 12940 17303
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 13280 16998 13308 17750
rect 13372 17134 13400 17818
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12728 14362 12756 16118
rect 12820 15706 12848 16458
rect 12912 15910 12940 16662
rect 13648 16425 13676 19654
rect 13740 18986 13768 20590
rect 14004 20392 14056 20398
rect 13910 20360 13966 20369
rect 14004 20334 14056 20340
rect 13910 20295 13966 20304
rect 13924 19718 13952 20295
rect 14016 20058 14044 20334
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13924 19310 13952 19654
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13924 19174 13952 19246
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13740 18958 13860 18986
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13740 18630 13768 18770
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13832 16969 13860 18958
rect 13924 18204 13952 19110
rect 14016 18358 14044 19994
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 13924 18176 14044 18204
rect 13818 16960 13874 16969
rect 13818 16895 13874 16904
rect 13634 16416 13690 16425
rect 13634 16351 13690 16360
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13358 15736 13414 15745
rect 12808 15700 12860 15706
rect 13358 15671 13360 15680
rect 12808 15642 12860 15648
rect 13412 15671 13414 15680
rect 13360 15642 13412 15648
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 15348 12940 15506
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 12820 15320 12940 15348
rect 12820 14482 12848 15320
rect 13082 15192 13138 15201
rect 13082 15127 13084 15136
rect 13136 15127 13138 15136
rect 13084 15098 13136 15104
rect 13280 15094 13308 15370
rect 13372 15366 13400 15642
rect 13648 15502 13676 15914
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13820 15632 13872 15638
rect 13740 15580 13820 15586
rect 13740 15574 13872 15580
rect 13740 15558 13860 15574
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13740 15008 13768 15558
rect 13648 14980 13768 15008
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12912 14362 12940 14418
rect 12728 14346 12940 14362
rect 12716 14340 12940 14346
rect 12768 14334 12940 14340
rect 12716 14282 12768 14288
rect 12728 13258 12756 14282
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 14074 13216 14214
rect 13556 14074 13584 14554
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12532 12436 12584 12442
rect 12820 12434 12848 13806
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13268 13388 13320 13394
rect 13320 13348 13400 13376
rect 13268 13330 13320 13336
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 12992 12776 13044 12782
rect 12990 12744 12992 12753
rect 13044 12744 13046 12753
rect 12990 12679 13046 12688
rect 13280 12646 13308 12786
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12532 12378 12584 12384
rect 12728 12406 12848 12434
rect 12530 12336 12586 12345
rect 12256 12300 12308 12306
rect 12530 12271 12586 12280
rect 12256 12242 12308 12248
rect 12268 12186 12296 12242
rect 12268 12158 12388 12186
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11898 12296 12038
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12268 10810 12296 11630
rect 12360 11218 12388 12158
rect 12544 11354 12572 12271
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 8634 12388 10542
rect 12452 9382 12480 10950
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8634 12572 8774
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12728 8514 12756 12406
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11286 12848 11834
rect 13280 11676 13308 12038
rect 13372 11830 13400 13348
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13280 11648 13400 11676
rect 13464 11665 13492 12038
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 13372 11218 13400 11648
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13464 11082 13492 11290
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10674 13492 11018
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13464 10198 13492 10610
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13556 10130 13584 13874
rect 13648 13802 13676 14980
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14618 13768 14826
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13924 13841 13952 15846
rect 13910 13832 13966 13841
rect 13636 13796 13688 13802
rect 13910 13767 13966 13776
rect 13636 13738 13688 13744
rect 14016 10470 14044 18176
rect 14108 17649 14136 21014
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14200 19718 14228 20946
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14200 19446 14228 19654
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14186 18728 14242 18737
rect 14186 18663 14242 18672
rect 14094 17640 14150 17649
rect 14094 17575 14150 17584
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14108 17338 14136 17478
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14108 12374 14136 17138
rect 14200 15450 14228 18663
rect 14292 17626 14320 23666
rect 14476 23225 14504 24142
rect 14462 23216 14518 23225
rect 14462 23151 14518 23160
rect 14370 23080 14426 23089
rect 14370 23015 14372 23024
rect 14424 23015 14426 23024
rect 14372 22986 14424 22992
rect 14476 22778 14504 23151
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14936 22094 14964 24958
rect 15028 22234 15056 26302
rect 15106 26200 15162 26302
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15106 23760 15162 23769
rect 15106 23695 15162 23704
rect 15120 23526 15148 23695
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 14936 22066 15056 22094
rect 15028 22030 15056 22066
rect 15396 22030 15424 24890
rect 15764 23798 15792 26200
rect 15844 25424 15896 25430
rect 15844 25366 15896 25372
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15488 22681 15516 23054
rect 15474 22672 15530 22681
rect 15474 22607 15530 22616
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14476 21010 14504 21354
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14476 20534 14504 20946
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14384 19718 14412 19926
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14370 19544 14426 19553
rect 14370 19479 14426 19488
rect 14384 19446 14412 19479
rect 14476 19446 14504 19790
rect 14568 19514 14596 19790
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14372 19236 14424 19242
rect 14372 19178 14424 19184
rect 14384 18902 14412 19178
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14476 18034 14504 19246
rect 14568 18358 14596 19450
rect 14660 18426 14688 20334
rect 15028 20058 15056 21286
rect 15120 21010 15148 21490
rect 15396 21457 15424 21558
rect 15382 21448 15438 21457
rect 15292 21412 15344 21418
rect 15382 21383 15438 21392
rect 15566 21448 15622 21457
rect 15566 21383 15568 21392
rect 15292 21354 15344 21360
rect 15620 21383 15622 21392
rect 15568 21354 15620 21360
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 19514 14872 19654
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15028 19310 15056 19994
rect 15304 19786 15332 21354
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15672 20806 15700 21286
rect 15660 20800 15712 20806
rect 15752 20800 15804 20806
rect 15660 20742 15712 20748
rect 15750 20768 15752 20777
rect 15804 20768 15806 20777
rect 15750 20703 15806 20712
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19922 15516 20198
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15106 19544 15162 19553
rect 15106 19479 15162 19488
rect 14832 19304 14884 19310
rect 14752 19264 14832 19292
rect 14752 18601 14780 19264
rect 14832 19246 14884 19252
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15120 19174 15148 19479
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14738 18592 14794 18601
rect 14738 18527 14794 18536
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14844 18358 14872 18906
rect 15016 18828 15068 18834
rect 15304 18816 15332 19722
rect 15856 19378 15884 25366
rect 15934 24712 15990 24721
rect 15934 24647 15990 24656
rect 15948 21690 15976 24647
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 17038 26330 17094 27000
rect 17682 26330 17738 27000
rect 17038 26302 17356 26330
rect 17038 26200 17094 26302
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 17144 24138 17172 24550
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 17132 24132 17184 24138
rect 17132 24074 17184 24080
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 17052 24018 17080 24074
rect 16960 23662 16988 24006
rect 17052 23990 17264 24018
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 16040 20466 16068 21082
rect 16132 20602 16160 22442
rect 16224 21486 16252 22442
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16224 20942 16252 21082
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16500 20505 16528 20810
rect 16486 20496 16542 20505
rect 16028 20460 16080 20466
rect 16486 20431 16542 20440
rect 16028 20402 16080 20408
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15068 18788 15332 18816
rect 15016 18770 15068 18776
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14832 18352 14884 18358
rect 14832 18294 14884 18300
rect 14936 18290 14964 18702
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15016 18624 15068 18630
rect 15014 18592 15016 18601
rect 15068 18592 15070 18601
rect 15014 18527 15070 18536
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15120 18329 15148 18362
rect 15106 18320 15162 18329
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 15016 18284 15068 18290
rect 15106 18255 15162 18264
rect 15016 18226 15068 18232
rect 14384 18006 14504 18034
rect 14554 18048 14610 18057
rect 14384 17814 14412 18006
rect 14554 17983 14610 17992
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14372 17808 14424 17814
rect 14476 17785 14504 17818
rect 14372 17750 14424 17756
rect 14462 17776 14518 17785
rect 14462 17711 14518 17720
rect 14292 17598 14412 17626
rect 14384 16794 14412 17598
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14370 16552 14426 16561
rect 14370 16487 14426 16496
rect 14384 16454 14412 16487
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14568 15450 14596 17983
rect 14936 17542 14964 18226
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14844 17082 14872 17478
rect 14752 17054 14872 17082
rect 14752 16114 14780 17054
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14200 15422 14412 15450
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14200 14822 14228 15302
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 14482 14228 14758
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14200 13258 14228 14418
rect 14292 14414 14320 14894
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 13326 14320 14350
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12442 14228 13194
rect 14292 12918 14320 13262
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14280 12776 14332 12782
rect 14384 12764 14412 15422
rect 14476 15422 14596 15450
rect 14476 14618 14504 15422
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14476 13802 14504 14554
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14332 12736 14412 12764
rect 14280 12718 14332 12724
rect 14292 12442 14320 12718
rect 14568 12646 14596 15302
rect 14660 13190 14688 16050
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14752 14929 14780 15030
rect 14738 14920 14794 14929
rect 14738 14855 14794 14864
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14200 11937 14228 12378
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14186 11928 14242 11937
rect 14186 11863 14242 11872
rect 14200 11830 14228 11863
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14200 11354 14228 11766
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14476 11150 14504 12106
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13832 9722 13860 10134
rect 14476 10062 14504 11086
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13648 9602 13676 9658
rect 13648 9574 13768 9602
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13360 8968 13412 8974
rect 13188 8916 13360 8922
rect 13188 8910 13412 8916
rect 13188 8906 13400 8910
rect 13176 8900 13400 8906
rect 13228 8894 13400 8900
rect 13176 8842 13228 8848
rect 12452 8486 12756 8514
rect 13556 8498 13584 9386
rect 13544 8492 13596 8498
rect 12452 8362 12480 8486
rect 13544 8434 13596 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12636 3466 12664 8366
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13372 7954 13400 8230
rect 13740 7954 13768 9574
rect 14476 9518 14504 9998
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8430 14596 9318
rect 14752 9110 14780 11698
rect 14844 10538 14872 16526
rect 14936 12850 14964 17478
rect 15028 17066 15056 18226
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15028 13530 15056 15506
rect 15120 15502 15148 15982
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15120 14618 15148 15030
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15120 13870 15148 14554
rect 15212 13938 15240 16594
rect 15396 16590 15424 17478
rect 15488 17134 15516 18634
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15382 16416 15438 16425
rect 15382 16351 15438 16360
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15094 15332 15914
rect 15396 15366 15424 16351
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15304 14822 15332 15030
rect 15292 14816 15344 14822
rect 15344 14776 15424 14804
rect 15292 14758 15344 14764
rect 15396 14346 15424 14776
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 13524 15068 13530
rect 15068 13484 15148 13512
rect 15016 13466 15068 13472
rect 15120 13002 15148 13484
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15028 12974 15148 13002
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14936 12714 14964 12786
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 12238 14964 12650
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15028 11694 15056 12974
rect 15212 12866 15240 13330
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15120 12838 15240 12866
rect 15120 12782 15148 12838
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15212 12306 15240 12718
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15198 11928 15254 11937
rect 15304 11914 15332 12582
rect 15396 12306 15424 12922
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15254 11886 15332 11914
rect 15198 11863 15200 11872
rect 15252 11863 15254 11872
rect 15200 11834 15252 11840
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 11082 15056 11494
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 15028 9926 15056 11018
rect 15212 11014 15240 11834
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15304 10810 15332 11494
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 10130 15240 10542
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15016 9920 15068 9926
rect 15304 9897 15332 9930
rect 15016 9862 15068 9868
rect 15290 9888 15346 9897
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 15028 8838 15056 9862
rect 15290 9823 15346 9832
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15396 8634 15424 10610
rect 15488 9110 15516 16934
rect 15580 16522 15608 18226
rect 16040 18086 16068 19314
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16224 19174 16252 19246
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16224 18086 16252 18634
rect 16408 18630 16436 19654
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16500 18902 16528 19178
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16486 18728 16542 18737
rect 16486 18663 16542 18672
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16500 18426 16528 18663
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15566 14784 15622 14793
rect 15566 14719 15622 14728
rect 15580 11898 15608 14719
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 10742 15700 17138
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15856 15638 15884 17070
rect 15948 15978 15976 17478
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 16040 15337 16068 18022
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16132 17338 16160 17682
rect 16224 17610 16252 18022
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16026 15328 16082 15337
rect 16026 15263 16082 15272
rect 16132 14958 16160 15846
rect 16120 14952 16172 14958
rect 15842 14920 15898 14929
rect 16120 14894 16172 14900
rect 15842 14855 15844 14864
rect 15896 14855 15898 14864
rect 15844 14826 15896 14832
rect 16316 14822 16344 16594
rect 16592 16590 16620 23190
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 21554 16712 22918
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16776 22438 16804 22578
rect 16868 22574 16896 23054
rect 16960 23050 16988 23598
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16762 21992 16818 22001
rect 16762 21927 16818 21936
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16776 21078 16804 21927
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16684 19242 16712 20742
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14482 16344 14758
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16500 14278 16528 16390
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 15094 16620 15302
rect 16684 15162 16712 16390
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16316 13258 16344 13670
rect 16408 13394 16436 14214
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16684 13734 16712 13942
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16684 12646 16712 13670
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16776 12434 16804 20198
rect 16868 18766 16896 22510
rect 17144 22234 17172 22646
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 16948 20800 17000 20806
rect 17052 20777 17080 21490
rect 16948 20742 17000 20748
rect 17038 20768 17094 20777
rect 16960 20602 16988 20742
rect 17038 20703 17094 20712
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17144 20330 17172 22170
rect 17236 20482 17264 23990
rect 17328 21486 17356 26302
rect 17420 26302 17738 26330
rect 17420 23186 17448 26302
rect 17682 26200 17738 26302
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26330 23534 27000
rect 24122 26330 24178 27000
rect 23478 26302 23704 26330
rect 23478 26200 23534 26302
rect 18144 24336 18196 24342
rect 17696 24284 18144 24290
rect 17696 24278 18196 24284
rect 17696 24262 18184 24278
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17406 22808 17462 22817
rect 17406 22743 17462 22752
rect 17420 22545 17448 22743
rect 17406 22536 17462 22545
rect 17406 22471 17462 22480
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17408 20936 17460 20942
rect 17406 20904 17408 20913
rect 17460 20904 17462 20913
rect 17406 20839 17462 20848
rect 17236 20454 17448 20482
rect 17512 20466 17540 21898
rect 17696 21690 17724 24262
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17972 23769 18000 23802
rect 18340 23798 18368 26200
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18328 23792 18380 23798
rect 17958 23760 18014 23769
rect 17958 23695 18014 23704
rect 18142 23760 18198 23769
rect 18328 23734 18380 23740
rect 18142 23695 18144 23704
rect 18196 23695 18198 23704
rect 18144 23666 18196 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17880 23322 17908 23598
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 18524 23118 18552 24074
rect 18708 23730 18736 24210
rect 18800 24070 18828 24550
rect 18984 24410 19012 26200
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18708 23526 18736 23666
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18524 22710 18552 23054
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17684 21412 17736 21418
rect 17684 21354 17736 21360
rect 17590 21312 17646 21321
rect 17590 21247 17646 21256
rect 17222 20360 17278 20369
rect 17132 20324 17184 20330
rect 17222 20295 17278 20304
rect 17132 20266 17184 20272
rect 17130 20088 17186 20097
rect 17236 20058 17264 20295
rect 17130 20023 17186 20032
rect 17224 20052 17276 20058
rect 16948 19712 17000 19718
rect 16946 19680 16948 19689
rect 17000 19680 17002 19689
rect 16946 19615 17002 19624
rect 17144 18873 17172 20023
rect 17224 19994 17276 20000
rect 17420 19836 17448 20454
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17604 20346 17632 21247
rect 17328 19808 17448 19836
rect 17512 20318 17632 20346
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17130 18864 17186 18873
rect 17130 18799 17186 18808
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18222 16988 18566
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16960 17746 16988 18158
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 17052 17218 17080 18158
rect 17144 17882 17172 18702
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17236 17746 17264 19110
rect 17328 17882 17356 19808
rect 17512 19666 17540 20318
rect 17420 19638 17540 19666
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17420 17626 17448 19638
rect 17500 19236 17552 19242
rect 17500 19178 17552 19184
rect 17512 18834 17540 19178
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17604 18290 17632 19654
rect 17696 19530 17724 21354
rect 17788 20806 17816 21626
rect 18432 21593 18460 22374
rect 18524 22166 18552 22646
rect 18800 22506 18828 24006
rect 19076 23798 19104 24278
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 19076 23254 19104 23734
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 18512 22160 18564 22166
rect 18512 22102 18564 22108
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 18524 22030 18552 22102
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18510 21720 18566 21729
rect 18510 21655 18566 21664
rect 18524 21622 18552 21655
rect 18512 21616 18564 21622
rect 18418 21584 18474 21593
rect 18512 21558 18564 21564
rect 18418 21519 18474 21528
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17776 20800 17828 20806
rect 17972 20788 18000 20946
rect 17776 20742 17828 20748
rect 17880 20760 18000 20788
rect 18328 20800 18380 20806
rect 17788 19990 17816 20742
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17774 19680 17830 19689
rect 17880 19666 17908 20760
rect 18328 20742 18380 20748
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 20262 18000 20334
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 18340 19854 18368 20742
rect 18418 20632 18474 20641
rect 18418 20567 18474 20576
rect 18432 20369 18460 20567
rect 18418 20360 18474 20369
rect 18418 20295 18474 20304
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 17830 19638 17908 19666
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18510 19680 18566 19689
rect 17774 19615 17830 19624
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17696 19502 17908 19530
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17880 19334 17908 19502
rect 18236 19372 18288 19378
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17696 19174 17724 19246
rect 17684 19168 17736 19174
rect 17682 19136 17684 19145
rect 17736 19136 17738 19145
rect 17682 19071 17738 19080
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 16960 17190 17080 17218
rect 17144 17598 17448 17626
rect 17144 17202 17172 17598
rect 17132 17196 17184 17202
rect 16960 16998 16988 17190
rect 17132 17138 17184 17144
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16868 14346 16896 15982
rect 16948 15904 17000 15910
rect 16946 15872 16948 15881
rect 17000 15872 17002 15881
rect 16946 15807 17002 15816
rect 17052 15570 17080 17002
rect 17236 16658 17264 17138
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17130 16280 17186 16289
rect 17130 16215 17186 16224
rect 17144 15910 17172 16215
rect 17328 15978 17356 16526
rect 17316 15972 17368 15978
rect 17316 15914 17368 15920
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17052 14464 17080 15506
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14929 17172 14962
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 17132 14476 17184 14482
rect 17052 14436 17132 14464
rect 17132 14418 17184 14424
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 17144 13938 17172 14418
rect 17236 14074 17264 14418
rect 17328 14074 17356 15370
rect 17420 15366 17448 17070
rect 17604 16114 17632 17750
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 14346 17448 15302
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16960 12986 16988 13874
rect 17144 13569 17172 13874
rect 17408 13864 17460 13870
rect 17512 13852 17540 15914
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17604 14890 17632 14962
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17460 13824 17540 13852
rect 17408 13806 17460 13812
rect 17130 13560 17186 13569
rect 17420 13530 17448 13806
rect 17498 13560 17554 13569
rect 17130 13495 17186 13504
rect 17408 13524 17460 13530
rect 17144 13394 17172 13495
rect 17498 13495 17554 13504
rect 17408 13466 17460 13472
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16592 12406 16804 12434
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11354 16160 11698
rect 16224 11354 16252 12242
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15764 9042 15792 10678
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16132 9382 16160 10542
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9722 16252 10066
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 16132 8922 16160 9318
rect 16132 8906 16252 8922
rect 16132 8900 16264 8906
rect 16132 8894 16212 8900
rect 16212 8842 16264 8848
rect 16316 8634 16344 10542
rect 16488 9920 16540 9926
rect 16486 9888 16488 9897
rect 16540 9888 16542 9897
rect 16486 9823 16542 9832
rect 16500 9654 16528 9823
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 8294 14780 8366
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 7546 13400 7686
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9416 800 9444 2450
rect 9784 2446 9812 2926
rect 10060 2854 10088 3062
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 11624 2582 11652 3334
rect 12820 3126 12848 5782
rect 14016 5778 14044 7142
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 15212 4146 15240 7958
rect 16592 7750 16620 12406
rect 17052 12306 17080 12582
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 12170 17080 12242
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11898 17448 12038
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10062 16896 11086
rect 17052 10810 17080 11630
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17328 10985 17356 11018
rect 17314 10976 17370 10985
rect 17314 10911 17370 10920
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16868 9518 16896 9998
rect 17052 9994 17080 10746
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 17328 9674 17356 10911
rect 17512 10674 17540 13495
rect 17604 11830 17632 14826
rect 17696 13852 17724 18022
rect 17788 15552 17816 19314
rect 17880 19310 18184 19334
rect 18236 19314 18288 19320
rect 17880 19306 18196 19310
rect 18144 19304 18196 19306
rect 18144 19246 18196 19252
rect 18052 19236 18104 19242
rect 18052 19178 18104 19184
rect 18064 18766 18092 19178
rect 18248 19145 18276 19314
rect 18234 19136 18290 19145
rect 18234 19071 18290 19080
rect 18340 18902 18368 19654
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17880 16114 17908 17274
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17788 15524 17908 15552
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17788 14822 17816 15370
rect 17880 14890 17908 15524
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17788 14328 17816 14758
rect 18340 14482 18368 16526
rect 18432 15162 18460 19654
rect 18510 19615 18566 19624
rect 18524 19514 18552 19615
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18510 18864 18566 18873
rect 18510 18799 18566 18808
rect 18524 18766 18552 18799
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 17134 18552 17478
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18524 16726 18552 17070
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18616 16590 18644 21286
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18708 18630 18736 20198
rect 18800 19174 18828 20946
rect 18892 20942 18920 21966
rect 19076 21486 19104 22102
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18892 20602 18920 20878
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18892 20398 18920 20538
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 18465 18736 18566
rect 18694 18456 18750 18465
rect 18694 18391 18750 18400
rect 18708 18057 18736 18391
rect 18694 18048 18750 18057
rect 18694 17983 18750 17992
rect 18800 17377 18828 18702
rect 18786 17368 18842 17377
rect 18786 17303 18842 17312
rect 18696 17264 18748 17270
rect 18748 17212 18828 17218
rect 18696 17206 18828 17212
rect 18708 17190 18828 17206
rect 18800 17134 18828 17190
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18892 16946 18920 20198
rect 18984 19922 19012 21422
rect 19062 21176 19118 21185
rect 19062 21111 19118 21120
rect 19076 20602 19104 21111
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18984 19378 19012 19722
rect 19076 19514 19104 19790
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18970 17368 19026 17377
rect 18970 17303 19026 17312
rect 18800 16918 18920 16946
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15434 18644 15846
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 17868 14340 17920 14346
rect 17788 14300 17868 14328
rect 17868 14282 17920 14288
rect 17880 14006 17908 14282
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17776 13864 17828 13870
rect 17696 13824 17776 13852
rect 17776 13806 17828 13812
rect 17880 13394 17908 13942
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 13258 17908 13330
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17774 13016 17830 13025
rect 17950 13019 18258 13028
rect 17774 12951 17830 12960
rect 17788 12753 17816 12951
rect 18340 12866 18368 13126
rect 18432 12918 18460 15098
rect 18800 14793 18828 16918
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18892 16046 18920 16730
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18880 14816 18932 14822
rect 18786 14784 18842 14793
rect 18880 14758 18932 14764
rect 18786 14719 18842 14728
rect 18892 14618 18920 14758
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18984 13818 19012 17303
rect 18616 13790 19012 13818
rect 18510 13560 18566 13569
rect 18510 13495 18566 13504
rect 18064 12838 18368 12866
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 17774 12744 17830 12753
rect 17774 12679 17830 12688
rect 17774 12608 17830 12617
rect 17774 12543 17830 12552
rect 17788 11898 17816 12543
rect 18064 12442 18092 12838
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18340 12170 18368 12242
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17144 9646 17356 9674
rect 17144 9518 17172 9646
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 16684 8838 16712 9454
rect 16868 9042 16896 9454
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15672 5234 15700 7210
rect 16868 5778 16896 8978
rect 17236 8090 17264 9454
rect 17604 8838 17632 11630
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17776 11008 17828 11014
rect 17774 10976 17776 10985
rect 17828 10976 17830 10985
rect 17774 10911 17830 10920
rect 17880 10742 17908 11018
rect 18432 11014 18460 12718
rect 18524 12714 18552 13495
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18616 12434 18644 13790
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12646 18736 12786
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18800 12442 18828 13398
rect 18984 13258 19012 13670
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18524 12406 18644 12434
rect 18788 12436 18840 12442
rect 18524 12102 18552 12406
rect 18788 12378 18840 12384
rect 18892 12170 18920 12854
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11626 18552 12038
rect 18602 11928 18658 11937
rect 18602 11863 18604 11872
rect 18656 11863 18658 11872
rect 18604 11834 18656 11840
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18984 11354 19012 13194
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18340 9450 18368 9862
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18432 8498 18460 9658
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18708 9382 18736 9590
rect 19076 9450 19104 19314
rect 19168 16114 19196 22374
rect 19260 20262 19288 22578
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19260 19514 19288 19858
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19260 14958 19288 17167
rect 19352 15450 19380 23598
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19444 22098 19472 22578
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19444 21350 19472 22034
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 20942 19472 21286
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19444 19281 19472 20402
rect 19430 19272 19486 19281
rect 19430 19207 19486 19216
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 18057 19472 18226
rect 19430 18048 19486 18057
rect 19430 17983 19486 17992
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19444 15570 19472 16526
rect 19536 16454 19564 24142
rect 19628 23322 19656 26200
rect 19982 24848 20038 24857
rect 19982 24783 20038 24792
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 19720 22778 19748 23258
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 20466 19656 21830
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 21010 19748 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 19922 19656 20266
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19720 19310 19748 19790
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18834 19748 19246
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19706 18728 19762 18737
rect 19706 18663 19762 18672
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 17610 19656 18158
rect 19616 17604 19668 17610
rect 19616 17546 19668 17552
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19628 15502 19656 15846
rect 19720 15745 19748 18663
rect 19706 15736 19762 15745
rect 19706 15671 19762 15680
rect 19616 15496 19668 15502
rect 19352 15422 19472 15450
rect 19616 15438 19668 15444
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19338 14920 19394 14929
rect 19338 14855 19394 14864
rect 19352 14822 19380 14855
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19168 12345 19196 12854
rect 19154 12336 19210 12345
rect 19154 12271 19210 12280
rect 19260 12186 19288 14418
rect 19168 12158 19288 12186
rect 19168 10198 19196 12158
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11150 19288 12038
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19168 9722 19196 10134
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 8838 18736 9318
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12084 800 12112 2450
rect 12452 2446 12480 2858
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14752 800 14780 2450
rect 15028 2446 15056 3878
rect 15488 3126 15516 5102
rect 16592 4826 16620 5578
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 16592 2854 16620 4762
rect 17052 3058 17080 5510
rect 17512 5234 17540 7142
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18708 5642 18736 8774
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17696 4486 17724 5102
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 3126 17724 4422
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17880 3058 17908 4966
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 19352 3466 19380 14758
rect 19444 14074 19472 15422
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19536 14822 19564 15030
rect 19720 15026 19748 15302
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19812 14906 19840 23054
rect 19904 20058 19932 24142
rect 19996 22094 20024 24783
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23186 20116 23462
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20088 22710 20116 23122
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 19996 22066 20116 22094
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19996 19786 20024 21898
rect 20088 21894 20116 22066
rect 20180 21978 20208 24346
rect 20272 22166 20300 26200
rect 20916 24274 20944 26200
rect 21270 24848 21326 24857
rect 21270 24783 21326 24792
rect 21086 24304 21142 24313
rect 20904 24268 20956 24274
rect 21086 24239 21142 24248
rect 20904 24210 20956 24216
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20364 22778 20392 22986
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20456 22094 20484 24006
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20548 22574 20576 23462
rect 20732 23032 20760 23734
rect 20812 23044 20864 23050
rect 20732 23004 20812 23032
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20640 22681 20668 22918
rect 20732 22710 20760 23004
rect 20812 22986 20864 22992
rect 20720 22704 20772 22710
rect 20626 22672 20682 22681
rect 20720 22646 20772 22652
rect 20626 22607 20682 22616
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20364 22066 20484 22094
rect 20364 22030 20392 22066
rect 20352 22024 20404 22030
rect 20180 21950 20300 21978
rect 20352 21966 20404 21972
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20166 21856 20222 21865
rect 20272 21842 20300 21950
rect 20272 21814 20484 21842
rect 20166 21791 20222 21800
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 15722 19932 19654
rect 20180 19530 20208 21791
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20272 21010 20300 21626
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20364 21321 20392 21422
rect 20350 21312 20406 21321
rect 20350 21247 20406 21256
rect 20260 21004 20312 21010
rect 20456 20992 20484 21814
rect 20260 20946 20312 20952
rect 20364 20964 20484 20992
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20272 19553 20300 19926
rect 20088 19502 20208 19530
rect 20258 19544 20314 19553
rect 20088 19446 20116 19502
rect 20258 19479 20314 19488
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19982 18592 20038 18601
rect 19982 18527 20038 18536
rect 19996 18222 20024 18527
rect 20088 18222 20116 18634
rect 20180 18358 20208 18838
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20272 18290 20300 18566
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19996 17785 20024 18158
rect 20074 17912 20130 17921
rect 20364 17898 20392 20964
rect 20640 20890 20668 22510
rect 21100 22094 21128 24239
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 21192 23866 21220 24142
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21100 22066 21220 22094
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20732 21350 20760 21558
rect 20812 21412 20864 21418
rect 20812 21354 20864 21360
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20456 20862 20668 20890
rect 20732 20874 20760 21286
rect 20720 20868 20772 20874
rect 20456 20806 20484 20862
rect 20720 20810 20772 20816
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 19922 20576 20742
rect 20732 20534 20760 20810
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20640 19310 20668 20334
rect 20732 19718 20760 20470
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 19446 20760 19654
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20074 17847 20130 17856
rect 20272 17870 20392 17898
rect 19982 17776 20038 17785
rect 19982 17711 20038 17720
rect 20088 16998 20116 17847
rect 20166 17640 20222 17649
rect 20166 17575 20222 17584
rect 20180 17270 20208 17575
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20272 15881 20300 17870
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20364 16658 20392 17682
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20456 16182 20484 17478
rect 20444 16176 20496 16182
rect 20444 16118 20496 16124
rect 20258 15872 20314 15881
rect 20258 15807 20314 15816
rect 19904 15694 20116 15722
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19720 14890 19840 14906
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19708 14884 19840 14890
rect 19760 14878 19840 14884
rect 19708 14826 19760 14832
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19628 14074 19656 14826
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19904 12374 19932 15370
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19892 12368 19944 12374
rect 19892 12310 19944 12316
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19720 11082 19748 11630
rect 19996 11218 20024 14962
rect 20088 13977 20116 15694
rect 20444 15360 20496 15366
rect 20548 15348 20576 18226
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17678 20668 18022
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20640 17066 20668 17478
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20732 16658 20760 17002
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20824 15910 20852 21354
rect 21192 20058 21220 22066
rect 21284 21729 21312 24783
rect 21362 24304 21418 24313
rect 21560 24274 21588 26200
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 21362 24239 21418 24248
rect 21548 24268 21600 24274
rect 21376 21962 21404 24239
rect 21548 24210 21600 24216
rect 22020 24206 22048 24754
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22112 23322 22140 24142
rect 22204 23497 22232 26200
rect 22848 25702 22876 26200
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22190 23488 22246 23497
rect 22190 23423 22246 23432
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22204 22778 22232 23258
rect 22296 23254 22324 23598
rect 22284 23248 22336 23254
rect 22284 23190 22336 23196
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22296 22642 22324 23054
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22572 22545 22600 24754
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22756 23032 22784 23734
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 23304 23336 23598
rect 23216 23276 23336 23304
rect 22836 23044 22888 23050
rect 22756 23004 22836 23032
rect 22836 22986 22888 22992
rect 23216 22692 23244 23276
rect 23308 23038 23520 23066
rect 23308 22982 23336 23038
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23400 22710 23428 22918
rect 23492 22710 23520 23038
rect 23676 22930 23704 26302
rect 24044 26302 24178 26330
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23584 22902 23704 22930
rect 23296 22704 23348 22710
rect 23216 22664 23296 22692
rect 23296 22646 23348 22652
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 22558 22536 22614 22545
rect 22558 22471 22614 22480
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21270 21720 21326 21729
rect 21270 21655 21326 21664
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20916 18272 20944 18634
rect 21008 18426 21036 19110
rect 21100 18902 21128 19110
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21468 18834 21496 19654
rect 21638 19544 21694 19553
rect 21638 19479 21694 19488
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21180 18284 21232 18290
rect 20916 18244 21180 18272
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20496 15337 20576 15348
rect 20496 15328 20590 15337
rect 20496 15320 20534 15328
rect 20444 15302 20496 15308
rect 20534 15263 20590 15272
rect 20640 15026 20668 15506
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20074 13968 20130 13977
rect 20074 13903 20130 13912
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 12986 20208 13670
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12306 20116 12718
rect 20364 12306 20392 13126
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10606 19748 11018
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10130 19748 10542
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19720 7818 19748 9930
rect 20180 9382 20208 10066
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20364 8430 20392 12242
rect 20456 8566 20484 13874
rect 20548 10470 20576 14214
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20732 12442 20760 13738
rect 20916 12753 20944 18244
rect 21180 18226 21232 18232
rect 21652 18170 21680 19479
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 21560 18142 21680 18170
rect 21008 17134 21036 18090
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 21100 17134 21128 17750
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21008 14006 21036 17070
rect 21100 16998 21128 17070
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21100 14618 21128 16934
rect 21192 16794 21220 17614
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21270 16144 21326 16153
rect 21270 16079 21326 16088
rect 21284 15910 21312 16079
rect 21376 15978 21404 16934
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21468 16250 21496 16458
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21560 16130 21588 18142
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21468 16102 21588 16130
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21100 14346 21128 14554
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21468 14278 21496 16102
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21192 12986 21220 14010
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21560 12850 21588 15846
rect 21652 15094 21680 16390
rect 21744 16046 21772 21830
rect 21836 21350 21864 22374
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21836 21078 21864 21286
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21836 18086 21864 21014
rect 22008 20528 22060 20534
rect 22112 20516 22140 21830
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22060 20488 22140 20516
rect 22008 20470 22060 20476
rect 22112 19242 22140 20488
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22020 18970 22048 19178
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21824 18080 21876 18086
rect 21928 18057 21956 18158
rect 21824 18022 21876 18028
rect 21914 18048 21970 18057
rect 21836 17882 21864 18022
rect 21914 17983 21970 17992
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21836 17202 21864 17818
rect 21928 17542 21956 17818
rect 22020 17814 22048 18770
rect 22112 18630 22140 19178
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 17270 21956 17478
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21836 16590 21864 17138
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21836 16266 21864 16526
rect 21836 16238 21956 16266
rect 21824 16176 21876 16182
rect 21822 16144 21824 16153
rect 21876 16144 21878 16153
rect 21822 16079 21878 16088
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21928 15638 21956 16238
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21652 13462 21680 13874
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21744 13326 21772 15574
rect 21928 15502 21956 15574
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14890 21956 15302
rect 22020 15026 22048 17614
rect 22112 15638 22140 18566
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 22112 15162 22140 15574
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21928 14346 21956 14826
rect 22020 14482 22048 14962
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 14006 21864 14214
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 21928 13530 21956 13670
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 22020 13326 22048 13874
rect 22204 13546 22232 20742
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22112 13518 22232 13546
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21744 12986 21772 13262
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21456 12776 21508 12782
rect 20902 12744 20958 12753
rect 21456 12718 21508 12724
rect 20902 12679 20958 12688
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20916 11898 20944 12582
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21468 11558 21496 12718
rect 21744 12170 21772 12922
rect 22112 12889 22140 13518
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22098 12880 22154 12889
rect 22204 12850 22232 13330
rect 22296 13297 22324 19654
rect 22282 13288 22338 13297
rect 22282 13223 22338 13232
rect 22098 12815 22154 12824
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12238 22232 12786
rect 22388 12434 22416 21830
rect 23308 21554 23336 22646
rect 23400 22574 23428 22646
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 21690 23520 22374
rect 23584 22137 23612 22902
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23570 22128 23626 22137
rect 23570 22063 23626 22072
rect 23676 21894 23704 22714
rect 23860 22094 23888 23462
rect 23940 22568 23992 22574
rect 24044 22545 24072 26302
rect 24122 26200 24178 26302
rect 24766 26200 24822 27000
rect 25410 26330 25466 27000
rect 25056 26302 25466 26330
rect 24214 24168 24270 24177
rect 24214 24103 24270 24112
rect 24490 24168 24546 24177
rect 24490 24103 24546 24112
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23940 22510 23992 22516
rect 24030 22536 24086 22545
rect 23768 22066 23888 22094
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22652 20800 22704 20806
rect 22756 20777 22784 20946
rect 22652 20742 22704 20748
rect 22742 20768 22798 20777
rect 22572 20262 22600 20742
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 22664 19446 22692 20742
rect 22742 20703 22798 20712
rect 23308 20466 23336 21490
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23400 20602 23428 20810
rect 23492 20806 23520 21286
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23676 20602 23704 20810
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22744 19372 22796 19378
rect 22744 19314 22796 19320
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22664 18970 22692 19246
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22480 18086 22508 18566
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 12714 22508 16390
rect 22572 13734 22600 17070
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22664 14958 22692 17002
rect 22756 16998 22784 19314
rect 22940 19174 22968 19926
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23308 19514 23336 19654
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 22928 19168 22980 19174
rect 22928 19110 22980 19116
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23400 18970 23428 19994
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23584 18766 23612 19450
rect 23676 18834 23704 19654
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 22834 18592 22890 18601
rect 22834 18527 22890 18536
rect 22848 18358 22876 18527
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22848 17338 22876 18294
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23584 17377 23612 17478
rect 23570 17368 23626 17377
rect 22836 17332 22888 17338
rect 23570 17303 23572 17312
rect 22836 17274 22888 17280
rect 23624 17303 23626 17312
rect 23572 17274 23624 17280
rect 23768 17252 23796 22066
rect 23952 21622 23980 22510
rect 24030 22471 24086 22480
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 24136 21146 24164 23054
rect 24228 21350 24256 24103
rect 24504 24070 24532 24103
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24400 23588 24452 23594
rect 24400 23530 24452 23536
rect 24412 23322 24440 23530
rect 24596 23526 24624 24006
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 24308 23316 24360 23322
rect 24308 23258 24360 23264
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24320 23186 24348 23258
rect 24780 23225 24808 26200
rect 25056 24274 25084 26302
rect 25410 26200 25466 26302
rect 26054 26330 26110 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 25780 24676 25832 24682
rect 25780 24618 25832 24624
rect 25964 24676 26016 24682
rect 25964 24618 26016 24624
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25148 24274 25176 24550
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25240 24138 25268 24210
rect 25320 24200 25372 24206
rect 25318 24168 25320 24177
rect 25372 24168 25374 24177
rect 25228 24132 25280 24138
rect 25318 24103 25374 24112
rect 25502 24168 25558 24177
rect 25502 24103 25558 24112
rect 25228 24074 25280 24080
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24964 23866 24992 24006
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 24766 23216 24822 23225
rect 24308 23180 24360 23186
rect 24766 23151 24822 23160
rect 24308 23122 24360 23128
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24398 22128 24454 22137
rect 24398 22063 24454 22072
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 19922 23888 20946
rect 24032 20800 24084 20806
rect 23952 20760 24032 20788
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23848 19440 23900 19446
rect 23848 19382 23900 19388
rect 23860 18970 23888 19382
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23846 18864 23902 18873
rect 23846 18799 23902 18808
rect 23676 17224 23796 17252
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22756 15094 22784 15302
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22664 13530 22692 14894
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22296 12406 22416 12434
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21744 11898 21772 12106
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10470 20668 10950
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 21192 9926 21220 11018
rect 21468 10810 21496 11494
rect 21744 11082 21772 11834
rect 22204 11694 22232 12174
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21744 10810 21772 11018
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21744 10198 21772 10746
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 9518 21220 9862
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 22204 7410 22232 11630
rect 22296 10266 22324 12406
rect 22756 11830 22784 14214
rect 22848 13870 22876 16594
rect 23308 16590 23336 16934
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 22926 16280 22982 16289
rect 22926 16215 22982 16224
rect 22940 16114 22968 16215
rect 23492 16182 23520 16390
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22848 11354 22876 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23112 13524 23164 13530
rect 23308 13512 23336 15438
rect 23584 15434 23612 16662
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23584 15162 23612 15370
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23164 13484 23336 13512
rect 23112 13466 23164 13472
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12986 22968 13126
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 23032 12850 23060 13262
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23584 12918 23612 13330
rect 23572 12912 23624 12918
rect 23572 12854 23624 12860
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22848 10606 22876 11290
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22572 7886 22600 9454
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23676 9081 23704 17224
rect 23860 16658 23888 18799
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23768 13462 23796 16390
rect 23860 15978 23888 16458
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23952 15706 23980 20760
rect 24032 20742 24084 20748
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24044 19786 24072 20334
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24044 18630 24072 18906
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 24044 18358 24072 18566
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 24044 17678 24072 18294
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24044 16250 24072 16526
rect 24136 16522 24164 19314
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24228 17785 24256 18566
rect 24214 17776 24270 17785
rect 24214 17711 24270 17720
rect 24228 17338 24256 17711
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23860 15162 23888 15302
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23860 14346 23888 15098
rect 23952 15026 23980 15370
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23952 14482 23980 14962
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23848 14340 23900 14346
rect 23900 14300 23980 14328
rect 23848 14282 23900 14288
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23860 13462 23888 13806
rect 23756 13456 23808 13462
rect 23756 13398 23808 13404
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23952 12918 23980 14300
rect 24044 13870 24072 15982
rect 24320 15910 24348 21286
rect 24412 21078 24440 22063
rect 24596 22001 24624 22918
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24688 22166 24716 22714
rect 24780 22642 24808 22986
rect 24952 22976 25004 22982
rect 25004 22936 25084 22964
rect 24952 22918 25004 22924
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 24582 21992 24638 22001
rect 24582 21927 24638 21936
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 21690 24624 21830
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 24780 21554 24808 22578
rect 24964 21876 24992 22578
rect 25056 22234 25084 22936
rect 25148 22710 25176 23598
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 25412 22500 25464 22506
rect 25412 22442 25464 22448
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 25056 21944 25084 22170
rect 25424 22030 25452 22442
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25228 21956 25280 21962
rect 25056 21916 25176 21944
rect 24964 21848 25084 21876
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24688 20398 24716 21422
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24780 20602 24808 20742
rect 25056 20618 25084 21848
rect 25148 21622 25176 21916
rect 25228 21898 25280 21904
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 25240 21554 25268 21898
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 24768 20596 24820 20602
rect 25056 20590 25268 20618
rect 24768 20538 24820 20544
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17746 24716 18022
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24398 17640 24454 17649
rect 24398 17575 24400 17584
rect 24452 17575 24454 17584
rect 24400 17546 24452 17552
rect 24596 17134 24624 17682
rect 24688 17202 24716 17682
rect 24872 17218 24900 19246
rect 24676 17196 24728 17202
rect 24872 17190 24992 17218
rect 24676 17138 24728 17144
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24688 17082 24716 17138
rect 24688 17054 24900 17082
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16182 24440 16934
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24504 15706 24532 16186
rect 24872 16114 24900 17054
rect 24964 16250 24992 17190
rect 25056 16590 25084 19654
rect 25148 18970 25176 20334
rect 25240 19786 25268 20590
rect 25318 20224 25374 20233
rect 25318 20159 25374 20168
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 16726 25176 17546
rect 25240 17542 25268 19722
rect 25332 19689 25360 20159
rect 25516 19854 25544 24103
rect 25792 24070 25820 24618
rect 25976 24138 26004 24618
rect 26068 24138 26096 24686
rect 26160 24313 26188 26302
rect 26698 26200 26754 27000
rect 27342 26330 27398 27000
rect 27986 26330 28042 27000
rect 27342 26302 27568 26330
rect 27342 26200 27398 26302
rect 26146 24304 26202 24313
rect 26146 24239 26202 24248
rect 26712 24138 26740 26200
rect 25964 24132 26016 24138
rect 25964 24074 26016 24080
rect 26056 24132 26108 24138
rect 26056 24074 26108 24080
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 27252 24064 27304 24070
rect 27252 24006 27304 24012
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25608 23050 25636 23734
rect 25688 23520 25740 23526
rect 25688 23462 25740 23468
rect 25596 23044 25648 23050
rect 25596 22986 25648 22992
rect 25700 22930 25728 23462
rect 26160 22982 26188 24006
rect 27172 23866 27200 24006
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 25608 22902 25728 22930
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 25608 22030 25636 22902
rect 25688 22772 25740 22778
rect 26252 22760 26280 23462
rect 27172 23186 27200 23598
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 26516 22976 26568 22982
rect 26516 22918 26568 22924
rect 25740 22732 26280 22760
rect 25688 22714 25740 22720
rect 26528 22438 26556 22918
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26528 22137 26556 22374
rect 27068 22160 27120 22166
rect 26514 22128 26570 22137
rect 26424 22092 26476 22098
rect 27068 22102 27120 22108
rect 26514 22063 26570 22072
rect 26424 22034 26476 22040
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25608 21010 25636 21966
rect 26436 21185 26464 22034
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26422 21176 26478 21185
rect 25976 21134 26372 21162
rect 25976 21078 26004 21134
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 25872 20800 25924 20806
rect 25686 20768 25742 20777
rect 25872 20742 25924 20748
rect 25686 20703 25742 20712
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25700 19786 25728 20703
rect 25884 20534 25912 20742
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 25318 19680 25374 19689
rect 25374 19638 25452 19666
rect 25318 19615 25374 19624
rect 25320 19236 25372 19242
rect 25320 19178 25372 19184
rect 25332 18358 25360 19178
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24308 15564 24360 15570
rect 24308 15506 24360 15512
rect 24320 14278 24348 15506
rect 24964 15162 24992 16186
rect 25056 16182 25084 16390
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 25134 16144 25190 16153
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25056 14906 25084 16118
rect 25134 16079 25190 16088
rect 25148 16046 25176 16079
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 25240 15570 25268 16594
rect 25332 16454 25360 16594
rect 25424 16454 25452 19638
rect 25700 18970 25728 19722
rect 25792 19310 25820 19790
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25870 19272 25926 19281
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25792 18834 25820 19246
rect 25870 19207 25926 19216
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25884 16658 25912 19207
rect 25976 18698 26004 20334
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 26068 18358 26096 20946
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26148 19916 26200 19922
rect 26148 19858 26200 19864
rect 26160 19258 26188 19858
rect 26252 19514 26280 20810
rect 26344 20330 26372 21134
rect 26422 21111 26478 21120
rect 26528 20856 26556 21898
rect 27080 21690 27108 22102
rect 27068 21684 27120 21690
rect 27068 21626 27120 21632
rect 26608 20868 26660 20874
rect 26528 20828 26608 20856
rect 26528 20466 26556 20828
rect 26608 20810 26660 20816
rect 27264 20602 27292 24006
rect 27540 23662 27568 26302
rect 27986 26302 28304 26330
rect 27986 26200 28042 26302
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27632 23186 27660 24278
rect 27712 23860 27764 23866
rect 27712 23802 27764 23808
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27724 23066 27752 23802
rect 27632 23038 27752 23066
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27356 22166 27384 22646
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27344 22160 27396 22166
rect 27448 22137 27476 22578
rect 27632 22574 27660 23038
rect 27710 22808 27766 22817
rect 27710 22743 27766 22752
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27724 22420 27752 22743
rect 27632 22392 27752 22420
rect 27344 22102 27396 22108
rect 27434 22128 27490 22137
rect 27434 22063 27490 22072
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 21690 27384 21830
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26332 20324 26384 20330
rect 26332 20266 26384 20272
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26344 19446 26372 20266
rect 26528 19768 26556 20402
rect 27448 20330 27476 22063
rect 27632 21078 27660 22392
rect 27816 22030 27844 25638
rect 28276 24682 28304 26302
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26330 29974 27000
rect 29918 26302 30144 26330
rect 29918 26200 29974 26302
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28644 24426 28672 26200
rect 29000 24608 29052 24614
rect 29092 24608 29144 24614
rect 29000 24550 29052 24556
rect 29090 24576 29092 24585
rect 29144 24576 29146 24585
rect 28644 24398 28856 24426
rect 28632 24268 28684 24274
rect 28632 24210 28684 24216
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 28184 23186 28212 23734
rect 28172 23180 28224 23186
rect 28172 23122 28224 23128
rect 28184 23050 28212 23122
rect 28172 23044 28224 23050
rect 28172 22986 28224 22992
rect 28368 22982 28396 24006
rect 28448 23588 28500 23594
rect 28448 23530 28500 23536
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 28460 22778 28488 23530
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28552 22710 28580 23190
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28644 22522 28672 24210
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28736 23322 28764 23462
rect 28724 23316 28776 23322
rect 28724 23258 28776 23264
rect 28736 22574 28764 23258
rect 28368 22494 28672 22522
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 28368 21894 28396 22494
rect 28448 22432 28500 22438
rect 28448 22374 28500 22380
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 28356 21548 28408 21554
rect 28460 21536 28488 22374
rect 28828 22234 28856 24398
rect 29012 23322 29040 24550
rect 29090 24511 29146 24520
rect 29182 24304 29238 24313
rect 29288 24274 29316 26200
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 29182 24239 29238 24248
rect 29276 24268 29328 24274
rect 29196 24206 29224 24239
rect 29276 24210 29328 24216
rect 30024 24206 30052 24754
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 29196 23526 29224 24142
rect 29552 24064 29604 24070
rect 29552 24006 29604 24012
rect 29564 23730 29592 24006
rect 30116 23798 30144 26302
rect 30562 26200 30618 27000
rect 31206 26330 31262 27000
rect 31206 26302 31340 26330
rect 31206 26200 31262 26302
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29184 23520 29236 23526
rect 29184 23462 29236 23468
rect 29552 23520 29604 23526
rect 29552 23462 29604 23468
rect 29000 23316 29052 23322
rect 29000 23258 29052 23264
rect 29092 23180 29144 23186
rect 29092 23122 29144 23128
rect 29104 22710 29132 23122
rect 29092 22704 29144 22710
rect 29092 22646 29144 22652
rect 29092 22432 29144 22438
rect 29092 22374 29144 22380
rect 28816 22228 28868 22234
rect 28816 22170 28868 22176
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28632 21888 28684 21894
rect 28632 21830 28684 21836
rect 28408 21508 28488 21536
rect 28356 21490 28408 21496
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27620 21072 27672 21078
rect 27620 21014 27672 21020
rect 27620 20936 27672 20942
rect 27540 20896 27620 20924
rect 27540 20641 27568 20896
rect 27620 20878 27672 20884
rect 27620 20800 27672 20806
rect 27908 20788 27936 21422
rect 27986 21176 28042 21185
rect 27986 21111 28042 21120
rect 28000 20806 28028 21111
rect 28092 20806 28120 21490
rect 28368 21010 28396 21490
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 27672 20760 27936 20788
rect 27988 20800 28040 20806
rect 27620 20742 27672 20748
rect 27988 20742 28040 20748
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 27526 20632 27582 20641
rect 27526 20567 27582 20576
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 26608 19780 26660 19786
rect 26528 19740 26608 19768
rect 26332 19440 26384 19446
rect 26332 19382 26384 19388
rect 26528 19378 26556 19740
rect 26608 19722 26660 19728
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26160 19230 26280 19258
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 26160 18465 26188 18770
rect 26146 18456 26202 18465
rect 26146 18391 26202 18400
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26160 16998 26188 18391
rect 26252 18222 26280 19230
rect 26240 18216 26292 18222
rect 26240 18158 26292 18164
rect 26252 17814 26280 18158
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26620 17105 26648 19450
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 26700 18896 26752 18902
rect 26700 18838 26752 18844
rect 26712 18601 26740 18838
rect 27172 18766 27200 19314
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 26698 18592 26754 18601
rect 26698 18527 26754 18536
rect 26804 18426 26832 18702
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26804 17610 26832 18362
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26804 17270 26832 17546
rect 26792 17264 26844 17270
rect 26792 17206 26844 17212
rect 26606 17096 26662 17105
rect 26606 17031 26662 17040
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 24872 14890 25084 14906
rect 24860 14884 25084 14890
rect 24912 14878 25084 14884
rect 24860 14826 24912 14832
rect 24964 14346 24992 14878
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 25044 14340 25096 14346
rect 25044 14282 25096 14288
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 23952 12646 23980 12854
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23952 12238 23980 12582
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 24044 12102 24072 13806
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11898 24072 12038
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23952 11354 23980 11766
rect 24136 11558 24164 13738
rect 24320 12782 24348 14214
rect 24596 14006 24624 14214
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24504 13258 24532 13466
rect 24492 13252 24544 13258
rect 24492 13194 24544 13200
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 12442 24440 12582
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24412 11898 24440 12378
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23952 9674 23980 11290
rect 24136 9994 24164 11494
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 23952 9646 24072 9674
rect 24596 9654 24624 13670
rect 25056 12170 25084 14282
rect 25240 13190 25268 15302
rect 25332 14346 25360 16390
rect 25424 16182 25452 16390
rect 26804 16250 26832 17206
rect 27080 16658 27108 18158
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 17610 27384 18022
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 27264 16658 27292 16934
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 15366 26096 15438
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 25596 15360 25648 15366
rect 25594 15328 25596 15337
rect 26056 15360 26108 15366
rect 25648 15328 25650 15337
rect 26056 15302 26108 15308
rect 25594 15263 25650 15272
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25332 14006 25360 14282
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25780 14272 25832 14278
rect 26068 14260 26096 15302
rect 26160 14414 26188 15370
rect 26804 15162 26832 16186
rect 27264 16046 27292 16594
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 26792 15156 26844 15162
rect 26792 15098 26844 15104
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14482 26648 14758
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26148 14272 26200 14278
rect 26068 14232 26148 14260
rect 25780 14214 25832 14220
rect 26148 14214 26200 14220
rect 25700 14006 25728 14214
rect 25792 14074 25820 14214
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25228 13184 25280 13190
rect 25228 13126 25280 13132
rect 26160 12753 26188 14214
rect 26146 12744 26202 12753
rect 26146 12679 26202 12688
rect 25044 12164 25096 12170
rect 25044 12106 25096 12112
rect 23662 9072 23718 9081
rect 23662 9007 23718 9016
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 5710 20944 6734
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 5778 22140 6598
rect 22480 5914 22508 7278
rect 22572 6322 22600 7822
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23952 7002 23980 7482
rect 24044 7478 24072 9646
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 24872 5778 24900 6054
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 20548 3058 20576 4966
rect 20916 4622 20944 5646
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5234 21404 5510
rect 22112 5234 22140 5714
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 27344 5636 27396 5642
rect 27344 5578 27396 5584
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 17420 800 17448 2450
rect 17512 2446 17540 2790
rect 20088 2446 20116 2790
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 1170 20208 2450
rect 22020 2446 22048 2790
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 25516 2650 25544 5578
rect 27172 5370 27200 5578
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 25976 4690 26004 4966
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 27356 2514 27384 5578
rect 27448 4672 27476 20266
rect 27632 19990 27660 20742
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27804 20528 27856 20534
rect 27710 20496 27766 20505
rect 27804 20470 27856 20476
rect 27710 20431 27766 20440
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27724 19922 27752 20431
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27540 19553 27568 19790
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27526 19544 27582 19553
rect 27526 19479 27582 19488
rect 27724 19378 27752 19654
rect 27712 19372 27764 19378
rect 27712 19314 27764 19320
rect 27816 19174 27844 20470
rect 28368 20466 28396 20946
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27620 18760 27672 18766
rect 27908 18714 27936 19246
rect 28368 19174 28396 19722
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 27620 18702 27672 18708
rect 27632 18329 27660 18702
rect 27816 18686 27936 18714
rect 27618 18320 27674 18329
rect 27816 18290 27844 18686
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27618 18255 27674 18264
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27526 17912 27582 17921
rect 27526 17847 27528 17856
rect 27580 17847 27582 17856
rect 27528 17818 27580 17824
rect 27816 17746 27844 18226
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27632 16250 27660 17478
rect 27816 17202 27844 17682
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27724 16590 27752 17070
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 27540 6798 27568 9522
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27540 5642 27568 6734
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27632 5574 27660 16186
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27816 7546 27844 11018
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 28368 5302 28396 19110
rect 28460 17898 28488 20878
rect 28552 20602 28580 21830
rect 28644 20913 28672 21830
rect 29012 21622 29040 21898
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 29104 21486 29132 22374
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 29196 21622 29224 21830
rect 29184 21616 29236 21622
rect 29184 21558 29236 21564
rect 29092 21480 29144 21486
rect 29092 21422 29144 21428
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28724 21072 28776 21078
rect 28724 21014 28776 21020
rect 28630 20904 28686 20913
rect 28630 20839 28686 20848
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28630 19952 28686 19961
rect 28630 19887 28632 19896
rect 28684 19887 28686 19896
rect 28632 19858 28684 19864
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28644 18358 28672 19110
rect 28736 18834 28764 21014
rect 28816 20800 28868 20806
rect 28816 20742 28868 20748
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 28632 18352 28684 18358
rect 28632 18294 28684 18300
rect 28460 17870 28580 17898
rect 28828 17882 28856 20742
rect 28920 20534 28948 21286
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28908 20528 28960 20534
rect 28908 20470 28960 20476
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28460 16522 28488 17750
rect 28552 16561 28580 17870
rect 28632 17876 28684 17882
rect 28632 17818 28684 17824
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28644 17218 28672 17818
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17338 28856 17478
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28644 17190 28856 17218
rect 28632 16720 28684 16726
rect 28632 16662 28684 16668
rect 28644 16590 28672 16662
rect 28632 16584 28684 16590
rect 28538 16552 28594 16561
rect 28448 16516 28500 16522
rect 28632 16526 28684 16532
rect 28538 16487 28594 16496
rect 28448 16458 28500 16464
rect 28644 16250 28672 16526
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 28828 12434 28856 17190
rect 28736 12406 28856 12434
rect 28736 6914 28764 12406
rect 28920 11121 28948 18702
rect 29012 16017 29040 20878
rect 29092 20528 29144 20534
rect 29196 20516 29224 21558
rect 29144 20488 29224 20516
rect 29092 20470 29144 20476
rect 29104 19718 29132 20470
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29104 19446 29132 19654
rect 29092 19440 29144 19446
rect 29092 19382 29144 19388
rect 29104 18970 29132 19382
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 29104 18358 29132 18906
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 29104 18170 29132 18294
rect 29104 18142 29224 18170
rect 29196 17746 29224 18142
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29196 17542 29224 17682
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29196 17202 29224 17478
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29564 16697 29592 23462
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 29736 22976 29788 22982
rect 29736 22918 29788 22924
rect 29748 19990 29776 22918
rect 30024 22506 30052 22986
rect 30012 22500 30064 22506
rect 30012 22442 30064 22448
rect 30024 21894 30052 22442
rect 30392 22438 30420 24686
rect 30576 24206 30604 26200
rect 31116 25016 31168 25022
rect 31116 24958 31168 24964
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 30932 24132 30984 24138
rect 30932 24074 30984 24080
rect 30944 23866 30972 24074
rect 31128 23866 31156 24958
rect 31208 24676 31260 24682
rect 31208 24618 31260 24624
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 31220 23730 31248 24618
rect 31208 23724 31260 23730
rect 31208 23666 31260 23672
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30484 23050 30512 23462
rect 30472 23044 30524 23050
rect 30472 22986 30524 22992
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 30472 21956 30524 21962
rect 30472 21898 30524 21904
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 30010 21584 30066 21593
rect 30010 21519 30066 21528
rect 30024 21010 30052 21519
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 30012 20392 30064 20398
rect 30300 20369 30328 21354
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30012 20334 30064 20340
rect 30286 20360 30342 20369
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29550 16688 29606 16697
rect 29550 16623 29606 16632
rect 28998 16008 29054 16017
rect 29748 15978 29776 18566
rect 29840 18086 29868 18702
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 28998 15943 29054 15952
rect 29736 15972 29788 15978
rect 29736 15914 29788 15920
rect 29932 15609 29960 19790
rect 30024 19174 30052 20334
rect 30286 20295 30342 20304
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30208 18834 30236 20198
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30300 19174 30328 19654
rect 30392 19514 30420 20742
rect 30484 19990 30512 21898
rect 30944 21554 30972 23598
rect 31220 23322 31248 23666
rect 31208 23316 31260 23322
rect 31208 23258 31260 23264
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31024 21888 31076 21894
rect 31024 21830 31076 21836
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30944 21350 30972 21490
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30668 21146 30696 21286
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30944 20874 30972 21286
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30472 19984 30524 19990
rect 30472 19926 30524 19932
rect 30484 19854 30512 19926
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30654 19408 30710 19417
rect 30654 19343 30656 19352
rect 30708 19343 30710 19352
rect 30656 19314 30708 19320
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30300 18970 30328 19110
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30116 18426 30144 18566
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30392 17814 30420 18090
rect 30668 17921 30696 18226
rect 30760 18222 30788 18634
rect 30840 18420 30892 18426
rect 30840 18362 30892 18368
rect 30852 18222 30880 18362
rect 30748 18216 30800 18222
rect 30748 18158 30800 18164
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30760 18086 30788 18158
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30654 17912 30710 17921
rect 30654 17847 30710 17856
rect 30380 17808 30432 17814
rect 30194 17776 30250 17785
rect 30380 17750 30432 17756
rect 30194 17711 30196 17720
rect 30248 17711 30250 17720
rect 30196 17682 30248 17688
rect 30102 17640 30158 17649
rect 30102 17575 30104 17584
rect 30156 17575 30158 17584
rect 30104 17546 30156 17552
rect 30116 17338 30144 17546
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 30208 17270 30236 17682
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30196 17264 30248 17270
rect 30196 17206 30248 17212
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30116 16998 30144 17138
rect 30300 16998 30328 17274
rect 30392 17134 30420 17750
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30852 17202 30880 17614
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30840 17196 30892 17202
rect 30840 17138 30892 17144
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30104 16992 30156 16998
rect 30104 16934 30156 16940
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 29918 15600 29974 15609
rect 29918 15535 29974 15544
rect 29736 13252 29788 13258
rect 29736 13194 29788 13200
rect 29748 11218 29776 13194
rect 30116 11354 30144 16934
rect 30852 16726 30880 17138
rect 30944 16794 30972 17478
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 30840 16720 30892 16726
rect 30840 16662 30892 16668
rect 31036 13433 31064 21830
rect 31114 21448 31170 21457
rect 31114 21383 31170 21392
rect 31128 20874 31156 21383
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 31220 17678 31248 22578
rect 31312 22506 31340 26302
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26330 33838 27000
rect 33782 26302 34100 26330
rect 33782 26200 33838 26302
rect 31576 25356 31628 25362
rect 31576 25298 31628 25304
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31392 24064 31444 24070
rect 31392 24006 31444 24012
rect 31300 22500 31352 22506
rect 31300 22442 31352 22448
rect 31300 21956 31352 21962
rect 31404 21944 31432 24006
rect 31496 23254 31524 24142
rect 31484 23248 31536 23254
rect 31484 23190 31536 23196
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31496 22778 31524 22918
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31496 22166 31524 22714
rect 31484 22160 31536 22166
rect 31484 22102 31536 22108
rect 31588 22098 31616 25298
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31668 22976 31720 22982
rect 31668 22918 31720 22924
rect 31680 22574 31708 22918
rect 31772 22778 31800 25094
rect 31864 24206 31892 26200
rect 32036 24880 32088 24886
rect 32036 24822 32088 24828
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 31864 23662 31892 24006
rect 31852 23656 31904 23662
rect 31852 23598 31904 23604
rect 32048 23322 32076 24822
rect 32508 24562 32536 26200
rect 32864 25560 32916 25566
rect 32864 25502 32916 25508
rect 32508 24534 32720 24562
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 32404 23656 32456 23662
rect 32126 23624 32182 23633
rect 32126 23559 32128 23568
rect 32180 23559 32182 23568
rect 32324 23616 32404 23644
rect 32128 23530 32180 23536
rect 32036 23316 32088 23322
rect 32036 23258 32088 23264
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31668 22568 31720 22574
rect 31668 22510 31720 22516
rect 31680 22166 31708 22510
rect 31668 22160 31720 22166
rect 31720 22108 31800 22114
rect 31668 22102 31800 22108
rect 31576 22092 31628 22098
rect 31680 22086 31800 22102
rect 32140 22094 32168 22986
rect 31576 22034 31628 22040
rect 31352 21916 31432 21944
rect 31300 21898 31352 21904
rect 31772 21554 31800 22086
rect 32048 22066 32168 22094
rect 32048 21894 32076 22066
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 32036 21888 32088 21894
rect 32036 21830 32088 21836
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 32048 21049 32076 21830
rect 32140 21418 32168 21966
rect 32128 21412 32180 21418
rect 32128 21354 32180 21360
rect 32034 21040 32090 21049
rect 32034 20975 32090 20984
rect 31760 20868 31812 20874
rect 31760 20810 31812 20816
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 31312 16658 31340 19858
rect 31772 19394 31800 20810
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31680 19366 31800 19394
rect 31680 18193 31708 19366
rect 31666 18184 31722 18193
rect 31666 18119 31722 18128
rect 31300 16652 31352 16658
rect 31300 16594 31352 16600
rect 31956 15473 31984 20742
rect 32324 19446 32352 23616
rect 32404 23598 32456 23604
rect 32508 22098 32536 24142
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32496 22092 32548 22098
rect 32496 22034 32548 22040
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32416 19825 32444 21490
rect 32496 21344 32548 21350
rect 32496 21286 32548 21292
rect 32402 19816 32458 19825
rect 32402 19751 32458 19760
rect 32312 19440 32364 19446
rect 32312 19382 32364 19388
rect 31942 15464 31998 15473
rect 31942 15399 31998 15408
rect 31022 13424 31078 13433
rect 32508 13394 32536 21286
rect 32600 21146 32628 23666
rect 32692 23322 32720 24534
rect 32876 23866 32904 25502
rect 33152 24664 33180 26200
rect 33600 25628 33652 25634
rect 33600 25570 33652 25576
rect 33506 24848 33562 24857
rect 33506 24783 33562 24792
rect 33152 24636 33364 24664
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33336 24206 33364 24636
rect 33520 24342 33548 24783
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32680 23316 32732 23322
rect 32680 23258 32732 23264
rect 33336 22778 33364 24142
rect 33612 23866 33640 25570
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33692 24948 33744 24954
rect 33692 24890 33744 24896
rect 33600 23860 33652 23866
rect 33600 23802 33652 23808
rect 33704 23118 33732 24890
rect 33796 23118 33824 25230
rect 34072 24342 34100 26302
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26330 37058 27000
rect 37002 26302 37228 26330
rect 37002 26200 37058 26302
rect 34244 25424 34296 25430
rect 34244 25366 34296 25372
rect 34060 24336 34112 24342
rect 34060 24278 34112 24284
rect 34072 24206 34100 24278
rect 34256 24274 34284 25366
rect 34440 24290 34468 26200
rect 34796 25220 34848 25226
rect 34796 25162 34848 25168
rect 34612 25084 34664 25090
rect 34612 25026 34664 25032
rect 34244 24268 34296 24274
rect 34440 24262 34560 24290
rect 34244 24210 34296 24216
rect 34532 24206 34560 24262
rect 34060 24200 34112 24206
rect 34060 24142 34112 24148
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34624 24070 34652 25026
rect 34612 24064 34664 24070
rect 34612 24006 34664 24012
rect 34808 23866 34836 25162
rect 35084 24206 35112 26200
rect 35624 25492 35676 25498
rect 35624 25434 35676 25440
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34980 23860 35032 23866
rect 34980 23802 35032 23808
rect 33874 23760 33930 23769
rect 33874 23695 33930 23704
rect 34888 23724 34940 23730
rect 33692 23112 33744 23118
rect 33692 23054 33744 23060
rect 33784 23112 33836 23118
rect 33784 23054 33836 23060
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 33324 22772 33376 22778
rect 33324 22714 33376 22720
rect 32954 22672 33010 22681
rect 32864 22636 32916 22642
rect 32954 22607 32956 22616
rect 32864 22578 32916 22584
rect 33008 22607 33010 22616
rect 32956 22578 33008 22584
rect 32876 22438 32904 22578
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32692 18902 32720 21354
rect 32680 18896 32732 18902
rect 32680 18838 32732 18844
rect 31022 13359 31078 13368
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 29736 11212 29788 11218
rect 29736 11154 29788 11160
rect 28906 11112 28962 11121
rect 30116 11082 30144 11290
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 28906 11047 28962 11056
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 31312 9654 31340 11086
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 32784 8401 32812 21966
rect 32876 9178 32904 22374
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 33336 18426 33364 22510
rect 33428 22438 33456 22986
rect 33888 22642 33916 23695
rect 34888 23666 34940 23672
rect 34612 23656 34664 23662
rect 34612 23598 34664 23604
rect 34428 23112 34480 23118
rect 34428 23054 34480 23060
rect 34518 23080 34574 23089
rect 34440 22794 34468 23054
rect 34518 23015 34574 23024
rect 34532 22982 34560 23015
rect 34520 22976 34572 22982
rect 34520 22918 34572 22924
rect 34440 22766 34560 22794
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 34532 22438 34560 22766
rect 33416 22432 33468 22438
rect 33416 22374 33468 22380
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 33324 18420 33376 18426
rect 33324 18362 33376 18368
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33428 15065 33456 22374
rect 34532 22234 34560 22374
rect 34520 22228 34572 22234
rect 34520 22170 34572 22176
rect 34624 19854 34652 23598
rect 34704 23588 34756 23594
rect 34704 23530 34756 23536
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34716 17678 34744 23530
rect 34900 22438 34928 23666
rect 34888 22432 34940 22438
rect 34888 22374 34940 22380
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 33414 15056 33470 15065
rect 33414 14991 33470 15000
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 34900 14618 34928 22374
rect 34992 20602 35020 23802
rect 35636 23798 35664 25434
rect 35728 24392 35756 26200
rect 35990 24712 36046 24721
rect 35900 24676 35952 24682
rect 35990 24647 36046 24656
rect 35900 24618 35952 24624
rect 35912 24392 35940 24618
rect 35728 24364 35940 24392
rect 35900 24132 35952 24138
rect 35900 24074 35952 24080
rect 35624 23792 35676 23798
rect 35624 23734 35676 23740
rect 35716 23112 35768 23118
rect 35716 23054 35768 23060
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35544 21690 35572 22918
rect 35728 22506 35756 23054
rect 35716 22500 35768 22506
rect 35716 22442 35768 22448
rect 35532 21684 35584 21690
rect 35532 21626 35584 21632
rect 34980 20596 35032 20602
rect 34980 20538 35032 20544
rect 35912 18737 35940 24074
rect 36004 23254 36032 24647
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 35992 23248 36044 23254
rect 35992 23190 36044 23196
rect 36004 23118 36032 23190
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 36096 22710 36124 23462
rect 36084 22704 36136 22710
rect 36084 22646 36136 22652
rect 36188 21962 36216 24006
rect 36372 23730 36400 26200
rect 36820 24676 36872 24682
rect 36820 24618 36872 24624
rect 36832 24206 36860 24618
rect 36820 24200 36872 24206
rect 37200 24188 37228 26302
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38934 26330 38990 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 37280 24200 37332 24206
rect 37200 24160 37280 24188
rect 36820 24142 36872 24148
rect 37280 24142 37332 24148
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36280 23322 36308 23666
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36268 23316 36320 23322
rect 36268 23258 36320 23264
rect 36176 21956 36228 21962
rect 36176 21898 36228 21904
rect 36544 21684 36596 21690
rect 36544 21626 36596 21632
rect 36556 21078 36584 21626
rect 36740 21622 36768 23462
rect 36832 23322 36860 24142
rect 37292 23322 37320 24142
rect 37464 24064 37516 24070
rect 37464 24006 37516 24012
rect 37476 23866 37504 24006
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37660 23730 37688 26200
rect 38488 24206 38516 26302
rect 38934 26302 39252 26330
rect 38934 26200 38990 26302
rect 39224 24206 39252 26302
rect 39578 26200 39634 27000
rect 40222 26330 40278 27000
rect 40866 26330 40922 27000
rect 40222 26302 40632 26330
rect 40222 26200 40278 26302
rect 39592 24274 39620 26200
rect 40316 24608 40368 24614
rect 40316 24550 40368 24556
rect 40328 24274 40356 24550
rect 39580 24268 39632 24274
rect 39580 24210 39632 24216
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 39212 24200 39264 24206
rect 39212 24142 39264 24148
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38488 23866 38516 24142
rect 39224 23866 39252 24142
rect 39304 24064 39356 24070
rect 39304 24006 39356 24012
rect 38476 23860 38528 23866
rect 38476 23802 38528 23808
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 36820 23316 36872 23322
rect 36820 23258 36872 23264
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 37832 23180 37884 23186
rect 37832 23122 37884 23128
rect 37844 22642 37872 23122
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37832 22636 37884 22642
rect 37832 22578 37884 22584
rect 39316 22001 39344 24006
rect 39592 23866 39620 24210
rect 40604 24206 40632 26302
rect 40866 26302 41184 26330
rect 40866 26200 40922 26302
rect 40592 24200 40644 24206
rect 40592 24142 40644 24148
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 39580 23860 39632 23866
rect 39580 23802 39632 23808
rect 40052 22778 40080 24074
rect 41156 23730 41184 26302
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 41524 24410 41552 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 41512 24404 41564 24410
rect 41512 24346 41564 24352
rect 41326 24168 41382 24177
rect 41326 24103 41382 24112
rect 41340 24070 41368 24103
rect 41328 24064 41380 24070
rect 41328 24006 41380 24012
rect 43456 23866 43484 26200
rect 43996 24064 44048 24070
rect 43996 24006 44048 24012
rect 43444 23860 43496 23866
rect 43444 23802 43496 23808
rect 41144 23724 41196 23730
rect 41144 23666 41196 23672
rect 41604 23656 41656 23662
rect 41604 23598 41656 23604
rect 41420 23520 41472 23526
rect 41420 23462 41472 23468
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40052 22234 40080 22714
rect 40040 22228 40092 22234
rect 40040 22170 40092 22176
rect 39302 21992 39358 22001
rect 39302 21927 39358 21936
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 36728 21616 36780 21622
rect 36728 21558 36780 21564
rect 36544 21072 36596 21078
rect 36544 21014 36596 21020
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 35898 18728 35954 18737
rect 35898 18663 35954 18672
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 41432 18086 41460 23462
rect 41616 18290 41644 23598
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 44008 18873 44036 24006
rect 44100 23746 44128 26200
rect 44744 24410 44772 26200
rect 44732 24404 44784 24410
rect 44732 24346 44784 24352
rect 44744 24206 44772 24346
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 46032 24206 46060 26200
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45284 24200 45336 24206
rect 45284 24142 45336 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 44100 23730 44220 23746
rect 44100 23724 44232 23730
rect 44100 23718 44180 23724
rect 44180 23666 44232 23672
rect 44456 23520 44508 23526
rect 44456 23462 44508 23468
rect 44468 19281 44496 23462
rect 44454 19272 44510 19281
rect 44454 19207 44510 19216
rect 43994 18864 44050 18873
rect 43994 18799 44050 18808
rect 41604 18284 41656 18290
rect 41604 18226 41656 18232
rect 41420 18080 41472 18086
rect 41420 18022 41472 18028
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 45296 17066 45324 24142
rect 45468 24064 45520 24070
rect 45468 24006 45520 24012
rect 45480 23662 45508 24006
rect 45572 23866 45600 24142
rect 45560 23860 45612 23866
rect 45560 23802 45612 23808
rect 46676 23730 46704 26200
rect 47320 24206 47348 26200
rect 47964 24206 47992 26200
rect 48318 24848 48374 24857
rect 48318 24783 48374 24792
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 47952 24200 48004 24206
rect 47952 24142 48004 24148
rect 46848 24064 46900 24070
rect 46848 24006 46900 24012
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 45468 23656 45520 23662
rect 45468 23598 45520 23604
rect 46860 20505 46888 24006
rect 47320 23866 47348 24142
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 48332 23730 48360 24783
rect 48320 23724 48372 23730
rect 48320 23666 48372 23672
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 48504 23520 48556 23526
rect 48504 23462 48556 23468
rect 46952 21690 46980 23462
rect 48412 22976 48464 22982
rect 48412 22918 48464 22924
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48424 22574 48452 22918
rect 48412 22568 48464 22574
rect 48412 22510 48464 22516
rect 48320 21888 48372 21894
rect 48320 21830 48372 21836
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 46940 21684 46992 21690
rect 46940 21626 46992 21632
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 47872 21350 47900 21490
rect 47860 21344 47912 21350
rect 47860 21286 47912 21292
rect 46846 20496 46902 20505
rect 46846 20431 46902 20440
rect 45284 17060 45336 17066
rect 45284 17002 45336 17008
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 34888 14612 34940 14618
rect 34888 14554 34940 14560
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 47872 11150 47900 21286
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48332 20058 48360 21830
rect 48516 21418 48544 23462
rect 48608 23118 48636 26200
rect 48688 24064 48740 24070
rect 48688 24006 48740 24012
rect 49516 24064 49568 24070
rect 49516 24006 49568 24012
rect 48596 23112 48648 23118
rect 48596 23054 48648 23060
rect 48608 22778 48636 23054
rect 48596 22772 48648 22778
rect 48596 22714 48648 22720
rect 48504 21412 48556 21418
rect 48504 21354 48556 21360
rect 48320 20052 48372 20058
rect 48320 19994 48372 20000
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 48700 15434 48728 24006
rect 49528 23905 49556 24006
rect 49514 23896 49570 23905
rect 49514 23831 49570 23840
rect 49528 23730 49556 23831
rect 49516 23724 49568 23730
rect 49516 23666 49568 23672
rect 49240 23520 49292 23526
rect 49240 23462 49292 23468
rect 48780 22976 48832 22982
rect 48780 22918 48832 22924
rect 48792 16998 48820 22918
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 48780 16992 48832 16998
rect 48780 16934 48832 16940
rect 48688 15428 48740 15434
rect 48688 15370 48740 15376
rect 49252 15366 49280 23462
rect 49332 23112 49384 23118
rect 49332 23054 49384 23060
rect 49344 22953 49372 23054
rect 49330 22944 49386 22953
rect 49330 22879 49386 22888
rect 49344 22778 49372 22879
rect 49332 22772 49384 22778
rect 49332 22714 49384 22720
rect 49516 22432 49568 22438
rect 49516 22374 49568 22380
rect 49528 22030 49556 22374
rect 49516 22024 49568 22030
rect 49514 21992 49516 22001
rect 49568 21992 49570 22001
rect 49514 21927 49570 21936
rect 49240 15360 49292 15366
rect 49240 15302 49292 15308
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47860 11144 47912 11150
rect 47860 11086 47912 11092
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 32864 9172 32916 9178
rect 32864 9114 32916 9120
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 32770 8392 32826 8401
rect 32770 8327 32826 8336
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 28736 6886 28948 6914
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 28356 5296 28408 5302
rect 28356 5238 28408 5244
rect 27528 4684 27580 4690
rect 27448 4644 27528 4672
rect 27528 4626 27580 4632
rect 27540 3602 27568 4626
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27816 2650 27844 4422
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 28552 3534 28580 5510
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28736 2650 28764 5714
rect 28920 5642 28948 6886
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 28908 5636 28960 5642
rect 28908 5578 28960 5584
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28828 4826 28856 5102
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28920 3670 28948 5578
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 41420 5160 41472 5166
rect 41420 5102 41472 5108
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33520 2650 33548 5034
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 27344 2508 27396 2514
rect 27344 2450 27396 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 20088 1142 20208 1170
rect 20088 800 20116 1142
rect 22756 800 22784 2450
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 25424 800 25452 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28092 870 28212 898
rect 28092 800 28120 870
rect 1398 0 1454 800
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 28184 762 28212 870
rect 28368 762 28396 2382
rect 30760 800 30788 2382
rect 33428 800 33456 2382
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 3402
rect 41432 800 41460 5102
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 44088 3664 44140 3670
rect 44088 3606 44140 3612
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 44100 800 44128 3606
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46768 800 46796 3538
rect 49424 3528 49476 3534
rect 49424 3470 49476 3476
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 3470
rect 28184 734 28396 762
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 1306 20712 1362 20768
rect 1398 19896 1454 19952
rect 1398 17856 1454 17912
rect 2778 24384 2834 24440
rect 1766 17312 1822 17368
rect 1214 17040 1270 17096
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1398 15272 1454 15328
rect 1306 15000 1362 15056
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 1306 13368 1362 13424
rect 1306 12180 1308 12200
rect 1308 12180 1360 12200
rect 1360 12180 1362 12200
rect 1306 12144 1362 12180
rect 1766 13932 1822 13968
rect 1766 13912 1768 13932
rect 1768 13912 1820 13932
rect 1820 13912 1822 13932
rect 1674 12552 1730 12608
rect 1582 11736 1638 11792
rect 1582 9696 1638 9752
rect 1766 8880 1822 8936
rect 2042 17448 2098 17504
rect 2042 16088 2098 16144
rect 3330 25608 3386 25664
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2686 21528 2742 21584
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3238 21936 3294 21992
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2686 19080 2742 19136
rect 2962 19488 3018 19544
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18672 2926 18728
rect 2778 18264 2834 18320
rect 2686 18128 2742 18184
rect 2594 14048 2650 14104
rect 2502 9288 2558 9344
rect 2410 8064 2466 8120
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2870 16632 2926 16688
rect 2778 13776 2834 13832
rect 4066 25200 4122 25256
rect 3606 24792 3662 24848
rect 3514 23976 3570 24032
rect 3514 22072 3570 22128
rect 3606 20576 3662 20632
rect 3606 20440 3662 20496
rect 3606 17876 3662 17912
rect 3606 17856 3608 17876
rect 3608 17856 3660 17876
rect 3660 17856 3662 17876
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 3514 14864 3570 14920
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3330 13252 3386 13288
rect 3330 13232 3332 13252
rect 3332 13232 3384 13252
rect 3384 13232 3386 13252
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 3330 11192 3386 11248
rect 2778 10920 2834 10976
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2870 10104 2926 10160
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2870 8472 2926 8528
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3606 12960 3662 13016
rect 4066 23588 4122 23624
rect 4066 23568 4068 23588
rect 4068 23568 4120 23588
rect 4120 23568 4122 23588
rect 4066 23160 4122 23216
rect 3882 22752 3938 22808
rect 3974 21120 4030 21176
rect 4158 22480 4214 22536
rect 4250 21004 4306 21040
rect 4250 20984 4252 21004
rect 4252 20984 4304 21004
rect 4304 20984 4306 21004
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 3606 11212 3662 11248
rect 3606 11192 3608 11212
rect 3608 11192 3660 11212
rect 3660 11192 3662 11212
rect 3606 10512 3662 10568
rect 3606 9560 3662 9616
rect 4066 15020 4122 15056
rect 4066 15000 4068 15020
rect 4068 15000 4120 15020
rect 4120 15000 4122 15020
rect 4434 17720 4490 17776
rect 4250 13504 4306 13560
rect 4158 12416 4214 12472
rect 4526 16496 4582 16552
rect 4434 15000 4490 15056
rect 4066 10004 4068 10024
rect 4068 10004 4120 10024
rect 4120 10004 4122 10024
rect 4066 9968 4122 10004
rect 4526 9560 4582 9616
rect 4710 16768 4766 16824
rect 5630 21548 5686 21584
rect 5630 21528 5632 21548
rect 5632 21528 5684 21548
rect 5684 21528 5686 21548
rect 5354 19352 5410 19408
rect 5354 17176 5410 17232
rect 5446 16632 5502 16688
rect 4710 13640 4766 13696
rect 5170 14592 5226 14648
rect 4986 11464 5042 11520
rect 4894 11328 4950 11384
rect 3698 7656 3754 7712
rect 2870 7248 2926 7304
rect 2778 6876 2780 6896
rect 2780 6876 2832 6896
rect 2832 6876 2834 6896
rect 2778 6840 2834 6876
rect 1306 6432 1362 6488
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 1306 6024 1362 6080
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 1306 5228 1362 5264
rect 1306 5208 1308 5228
rect 1308 5208 1360 5228
rect 1360 5208 1362 5228
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 1306 4800 1362 4856
rect 1766 4392 1822 4448
rect 3514 4392 3570 4448
rect 2686 4120 2742 4176
rect 2870 3984 2926 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 3576 1362 3632
rect 1306 3168 1362 3224
rect 1306 2760 1362 2816
rect 1306 2352 1362 2408
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2778 1944 2834 2000
rect 3330 1536 3386 1592
rect 5630 19896 5686 19952
rect 5630 17856 5686 17912
rect 6550 24112 6606 24168
rect 6182 21528 6238 21584
rect 6734 23468 6736 23488
rect 6736 23468 6788 23488
rect 6788 23468 6790 23488
rect 6734 23432 6790 23468
rect 6274 20712 6330 20768
rect 5906 17076 5908 17096
rect 5908 17076 5960 17096
rect 5960 17076 5962 17096
rect 5906 17040 5962 17076
rect 5722 15816 5778 15872
rect 5538 14728 5594 14784
rect 5354 10512 5410 10568
rect 5722 14456 5778 14512
rect 6642 22072 6698 22128
rect 6550 19896 6606 19952
rect 6458 19372 6514 19408
rect 6458 19352 6460 19372
rect 6460 19352 6512 19372
rect 6512 19352 6514 19372
rect 6274 17856 6330 17912
rect 6090 16496 6146 16552
rect 6550 17584 6606 17640
rect 6458 17312 6514 17368
rect 6550 17040 6606 17096
rect 6458 16632 6514 16688
rect 6182 15020 6238 15056
rect 6182 15000 6184 15020
rect 6184 15000 6236 15020
rect 6236 15000 6238 15020
rect 7194 23568 7250 23624
rect 6918 19216 6974 19272
rect 6734 16496 6790 16552
rect 6550 15816 6606 15872
rect 6642 15544 6698 15600
rect 6182 11056 6238 11112
rect 6366 10376 6422 10432
rect 7194 17992 7250 18048
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8114 20848 8170 20904
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 9126 24792 9182 24848
rect 8666 21528 8722 21584
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7470 16496 7526 16552
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7194 15444 7196 15464
rect 7196 15444 7248 15464
rect 7248 15444 7250 15464
rect 7194 15408 7250 15444
rect 7102 12824 7158 12880
rect 7010 11464 7066 11520
rect 7562 15680 7618 15736
rect 7194 12552 7250 12608
rect 7654 15272 7710 15328
rect 8022 16788 8078 16824
rect 8022 16768 8024 16788
rect 8024 16768 8076 16788
rect 8076 16768 8078 16788
rect 8114 16632 8170 16688
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8390 16088 8446 16144
rect 8482 15952 8538 16008
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7654 14900 7656 14920
rect 7656 14900 7708 14920
rect 7708 14900 7710 14920
rect 7654 14864 7710 14900
rect 7838 15000 7894 15056
rect 7286 10648 7342 10704
rect 7194 9172 7250 9208
rect 7194 9152 7196 9172
rect 7196 9152 7248 9172
rect 7248 9152 7250 9172
rect 6274 4140 6330 4176
rect 6274 4120 6276 4140
rect 6276 4120 6328 4140
rect 6328 4120 6330 4140
rect 7746 12552 7802 12608
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 8206 11772 8208 11792
rect 8208 11772 8260 11792
rect 8260 11772 8262 11792
rect 8206 11736 8262 11772
rect 8666 15544 8722 15600
rect 9218 17992 9274 18048
rect 9034 17040 9090 17096
rect 8758 14728 8814 14784
rect 8574 14592 8630 14648
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7746 9016 7802 9072
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 8758 11736 8814 11792
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 9218 15564 9274 15600
rect 9218 15544 9220 15564
rect 9220 15544 9272 15564
rect 9272 15544 9274 15564
rect 9770 21292 9772 21312
rect 9772 21292 9824 21312
rect 9824 21292 9826 21312
rect 9770 21256 9826 21292
rect 9402 20440 9458 20496
rect 10230 21412 10286 21448
rect 10230 21392 10232 21412
rect 10232 21392 10284 21412
rect 10284 21392 10286 21412
rect 9494 18400 9550 18456
rect 9586 17856 9642 17912
rect 9494 15680 9550 15736
rect 9494 14456 9550 14512
rect 9770 18808 9826 18864
rect 9954 17312 10010 17368
rect 9770 17176 9826 17232
rect 9678 15816 9734 15872
rect 10414 19352 10470 19408
rect 11886 24248 11942 24304
rect 11886 23468 11888 23488
rect 11888 23468 11940 23488
rect 11940 23468 11942 23488
rect 11886 23432 11942 23468
rect 11794 22752 11850 22808
rect 11242 21392 11298 21448
rect 10046 16088 10102 16144
rect 9862 15952 9918 16008
rect 9862 15428 9918 15464
rect 9862 15408 9864 15428
rect 9864 15408 9916 15428
rect 9916 15408 9918 15428
rect 9862 15136 9918 15192
rect 9494 13504 9550 13560
rect 9402 13388 9458 13424
rect 9402 13368 9404 13388
rect 9404 13368 9456 13388
rect 9456 13368 9458 13388
rect 10046 14764 10048 14784
rect 10048 14764 10100 14784
rect 10100 14764 10102 14784
rect 10046 14728 10102 14764
rect 10322 16088 10378 16144
rect 9770 11600 9826 11656
rect 9770 11328 9826 11384
rect 9310 11056 9366 11112
rect 9586 8356 9642 8392
rect 9586 8336 9588 8356
rect 9588 8336 9640 8356
rect 9640 8336 9642 8356
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 10966 18672 11022 18728
rect 10874 18536 10930 18592
rect 11334 20712 11390 20768
rect 11058 17176 11114 17232
rect 11150 16904 11206 16960
rect 11058 16496 11114 16552
rect 10874 16088 10930 16144
rect 10966 15972 11022 16008
rect 10966 15952 10968 15972
rect 10968 15952 11020 15972
rect 11020 15952 11022 15972
rect 11058 15272 11114 15328
rect 10966 15136 11022 15192
rect 10782 13776 10838 13832
rect 10690 12844 10746 12880
rect 10690 12824 10692 12844
rect 10692 12824 10744 12844
rect 10744 12824 10746 12844
rect 10230 10920 10286 10976
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 11334 14900 11336 14920
rect 11336 14900 11388 14920
rect 11388 14900 11390 14920
rect 11334 14864 11390 14900
rect 11794 19760 11850 19816
rect 12254 23568 12310 23624
rect 11886 18400 11942 18456
rect 11058 11192 11114 11248
rect 11610 12960 11666 13016
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13910 21120 13966 21176
rect 12346 18672 12402 18728
rect 13358 20168 13414 20224
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12438 18264 12494 18320
rect 12162 18128 12218 18184
rect 12070 17584 12126 17640
rect 12438 16632 12494 16688
rect 12070 16224 12126 16280
rect 12070 15580 12072 15600
rect 12072 15580 12124 15600
rect 12124 15580 12126 15600
rect 12070 15544 12126 15580
rect 11978 15020 12034 15056
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 12070 14728 12126 14784
rect 11978 11736 12034 11792
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13634 20304 13690 20360
rect 13634 20032 13690 20088
rect 13542 17856 13598 17912
rect 12898 17312 12954 17368
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13910 20304 13966 20360
rect 13818 16904 13874 16960
rect 13634 16360 13690 16416
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13358 15700 13414 15736
rect 13358 15680 13360 15700
rect 13360 15680 13412 15700
rect 13412 15680 13414 15700
rect 13082 15156 13138 15192
rect 13082 15136 13084 15156
rect 13084 15136 13136 15156
rect 13136 15136 13138 15156
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12990 12724 12992 12744
rect 12992 12724 13044 12744
rect 13044 12724 13046 12744
rect 12990 12688 13046 12724
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12530 12280 12586 12336
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13450 11600 13506 11656
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13910 13776 13966 13832
rect 14186 18672 14242 18728
rect 14094 17584 14150 17640
rect 14462 23160 14518 23216
rect 14370 23044 14426 23080
rect 14370 23024 14372 23044
rect 14372 23024 14424 23044
rect 14424 23024 14426 23044
rect 15106 23704 15162 23760
rect 15474 22616 15530 22672
rect 14370 19488 14426 19544
rect 15382 21392 15438 21448
rect 15566 21412 15622 21448
rect 15566 21392 15568 21412
rect 15568 21392 15620 21412
rect 15620 21392 15622 21412
rect 15750 20748 15752 20768
rect 15752 20748 15804 20768
rect 15804 20748 15806 20768
rect 15750 20712 15806 20748
rect 15106 19488 15162 19544
rect 14738 18536 14794 18592
rect 15934 24656 15990 24712
rect 16486 20440 16542 20496
rect 15014 18572 15016 18592
rect 15016 18572 15068 18592
rect 15068 18572 15070 18592
rect 15014 18536 15070 18572
rect 15106 18264 15162 18320
rect 14554 17992 14610 18048
rect 14462 17720 14518 17776
rect 14370 16496 14426 16552
rect 14738 14864 14794 14920
rect 14186 11872 14242 11928
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 15382 16360 15438 16416
rect 15198 11892 15254 11928
rect 15198 11872 15200 11892
rect 15200 11872 15252 11892
rect 15252 11872 15254 11892
rect 15290 9832 15346 9888
rect 16486 18672 16542 18728
rect 15566 14728 15622 14784
rect 16026 15272 16082 15328
rect 15842 14884 15898 14920
rect 15842 14864 15844 14884
rect 15844 14864 15896 14884
rect 15896 14864 15898 14884
rect 16762 21936 16818 21992
rect 17038 20712 17094 20768
rect 17406 22752 17462 22808
rect 17406 22480 17462 22536
rect 17406 20884 17408 20904
rect 17408 20884 17460 20904
rect 17460 20884 17462 20904
rect 17406 20848 17462 20884
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17958 23704 18014 23760
rect 18142 23724 18198 23760
rect 18142 23704 18144 23724
rect 18144 23704 18196 23724
rect 18196 23704 18198 23724
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17590 21256 17646 21312
rect 17222 20304 17278 20360
rect 17130 20032 17186 20088
rect 16946 19660 16948 19680
rect 16948 19660 17000 19680
rect 17000 19660 17002 19680
rect 16946 19624 17002 19660
rect 17130 18808 17186 18864
rect 18510 21664 18566 21720
rect 18418 21528 18474 21584
rect 17774 19624 17830 19680
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18418 20576 18474 20632
rect 18418 20304 18474 20360
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17682 19116 17684 19136
rect 17684 19116 17736 19136
rect 17736 19116 17738 19136
rect 17682 19080 17738 19116
rect 16946 15852 16948 15872
rect 16948 15852 17000 15872
rect 17000 15852 17002 15872
rect 16946 15816 17002 15852
rect 17130 16224 17186 16280
rect 17130 14864 17186 14920
rect 17130 13504 17186 13560
rect 17498 13504 17554 13560
rect 16486 9868 16488 9888
rect 16488 9868 16540 9888
rect 16540 9868 16542 9888
rect 16486 9832 16542 9868
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 17314 10920 17370 10976
rect 18234 19080 18290 19136
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18510 19624 18566 19680
rect 18510 18808 18566 18864
rect 18694 18400 18750 18456
rect 18694 17992 18750 18048
rect 18786 17312 18842 17368
rect 19062 21120 19118 21176
rect 18970 17312 19026 17368
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17774 12960 17830 13016
rect 18786 14728 18842 14784
rect 18510 13504 18566 13560
rect 17774 12688 17830 12744
rect 17774 12552 17830 12608
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17774 10956 17776 10976
rect 17776 10956 17828 10976
rect 17828 10956 17830 10976
rect 17774 10920 17830 10956
rect 18602 11892 18658 11928
rect 18602 11872 18604 11892
rect 18604 11872 18656 11892
rect 18656 11872 18658 11892
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 19246 17176 19302 17232
rect 19430 19216 19486 19272
rect 19430 17992 19486 18048
rect 19982 24792 20038 24848
rect 19706 18672 19762 18728
rect 19706 15680 19762 15736
rect 19338 14864 19394 14920
rect 19154 12280 19210 12336
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 21270 24792 21326 24848
rect 21086 24248 21142 24304
rect 20626 22616 20682 22672
rect 20166 21800 20222 21856
rect 20350 21256 20406 21312
rect 20258 19488 20314 19544
rect 19982 18536 20038 18592
rect 20074 17856 20130 17912
rect 19982 17720 20038 17776
rect 20166 17584 20222 17640
rect 20258 15816 20314 15872
rect 21362 24248 21418 24304
rect 22190 23432 22246 23488
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22558 22480 22614 22536
rect 21270 21664 21326 21720
rect 21638 19488 21694 19544
rect 20534 15272 20590 15328
rect 20074 13912 20130 13968
rect 21270 16088 21326 16144
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 21914 17992 21970 18048
rect 21822 16124 21824 16144
rect 21824 16124 21876 16144
rect 21876 16124 21878 16144
rect 21822 16088 21878 16124
rect 20902 12688 20958 12744
rect 22098 12824 22154 12880
rect 22282 13232 22338 13288
rect 23570 22072 23626 22128
rect 24214 24112 24270 24168
rect 24490 24112 24546 24168
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22742 20712 22798 20768
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22834 18536 22890 18592
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23570 17332 23626 17368
rect 23570 17312 23572 17332
rect 23572 17312 23624 17332
rect 23624 17312 23626 17332
rect 24030 22480 24086 22536
rect 25318 24148 25320 24168
rect 25320 24148 25372 24168
rect 25372 24148 25374 24168
rect 25318 24112 25374 24148
rect 25502 24112 25558 24168
rect 24766 23160 24822 23216
rect 24398 22072 24454 22128
rect 23846 18808 23902 18864
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22926 16224 22982 16280
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 24214 17720 24270 17776
rect 24582 21936 24638 21992
rect 24398 17604 24454 17640
rect 24398 17584 24400 17604
rect 24400 17584 24452 17604
rect 24452 17584 24454 17604
rect 25318 20168 25374 20224
rect 26146 24248 26202 24304
rect 26514 22072 26570 22128
rect 25686 20712 25742 20768
rect 25318 19624 25374 19680
rect 25134 16088 25190 16144
rect 25870 19216 25926 19272
rect 26422 21120 26478 21176
rect 27710 22752 27766 22808
rect 27434 22072 27490 22128
rect 29090 24556 29092 24576
rect 29092 24556 29144 24576
rect 29144 24556 29146 24576
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 29090 24520 29146 24556
rect 29182 24248 29238 24304
rect 27986 21120 28042 21176
rect 27526 20576 27582 20632
rect 26146 18400 26202 18456
rect 26698 18536 26754 18592
rect 26606 17040 26662 17096
rect 25594 15308 25596 15328
rect 25596 15308 25648 15328
rect 25648 15308 25650 15328
rect 25594 15272 25650 15308
rect 26146 12688 26202 12744
rect 23662 9016 23718 9072
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27710 20440 27766 20496
rect 27526 19488 27582 19544
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27618 18264 27674 18320
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27526 17876 27582 17912
rect 27526 17856 27528 17876
rect 27528 17856 27580 17876
rect 27580 17856 27582 17876
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 28630 20848 28686 20904
rect 28630 19916 28686 19952
rect 28630 19896 28632 19916
rect 28632 19896 28684 19916
rect 28684 19896 28686 19916
rect 28538 16496 28594 16552
rect 30010 21528 30066 21584
rect 29550 16632 29606 16688
rect 28998 15952 29054 16008
rect 30286 20304 30342 20360
rect 30654 19372 30710 19408
rect 30654 19352 30656 19372
rect 30656 19352 30708 19372
rect 30708 19352 30710 19372
rect 30654 17856 30710 17912
rect 30194 17740 30250 17776
rect 30194 17720 30196 17740
rect 30196 17720 30248 17740
rect 30248 17720 30250 17740
rect 30102 17604 30158 17640
rect 30102 17584 30104 17604
rect 30104 17584 30156 17604
rect 30156 17584 30158 17604
rect 29918 15544 29974 15600
rect 31114 21392 31170 21448
rect 32126 23588 32182 23624
rect 32126 23568 32128 23588
rect 32128 23568 32180 23588
rect 32180 23568 32182 23588
rect 32034 20984 32090 21040
rect 31666 18128 31722 18184
rect 32402 19760 32458 19816
rect 31942 15408 31998 15464
rect 31022 13368 31078 13424
rect 33506 24792 33562 24848
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33874 23704 33930 23760
rect 32954 22636 33010 22672
rect 32954 22616 32956 22636
rect 32956 22616 33008 22636
rect 33008 22616 33010 22636
rect 28906 11056 28962 11112
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 34518 23024 34574 23080
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 33414 15000 33470 15056
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 35990 24656 36046 24712
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 41326 24112 41382 24168
rect 39302 21936 39358 21992
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 35898 18672 35954 18728
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 44454 19216 44510 19272
rect 43994 18808 44050 18864
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 48318 24792 48374 24848
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 46846 20440 46902 20496
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49514 23840 49570 23896
rect 49146 20984 49202 21040
rect 49330 22888 49386 22944
rect 49514 21972 49516 21992
rect 49516 21972 49568 21992
rect 49568 21972 49570 21992
rect 49514 21936 49570 21972
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 32770 8336 32826 8392
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3325 25666 3391 25669
rect 0 25664 3391 25666
rect 0 25608 3330 25664
rect 3386 25608 3391 25664
rect 0 25606 3391 25608
rect 0 25576 800 25606
rect 3325 25603 3391 25606
rect 0 25258 800 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 800 25198
rect 4061 25195 4127 25198
rect 0 24850 800 24880
rect 3601 24850 3667 24853
rect 0 24848 3667 24850
rect 0 24792 3606 24848
rect 3662 24792 3667 24848
rect 0 24790 3667 24792
rect 0 24760 800 24790
rect 3601 24787 3667 24790
rect 9121 24850 9187 24853
rect 19977 24850 20043 24853
rect 9121 24848 20043 24850
rect 9121 24792 9126 24848
rect 9182 24792 19982 24848
rect 20038 24792 20043 24848
rect 9121 24790 20043 24792
rect 9121 24787 9187 24790
rect 19977 24787 20043 24790
rect 21265 24850 21331 24853
rect 33501 24850 33567 24853
rect 21265 24848 33567 24850
rect 21265 24792 21270 24848
rect 21326 24792 33506 24848
rect 33562 24792 33567 24848
rect 21265 24790 33567 24792
rect 21265 24787 21331 24790
rect 33501 24787 33567 24790
rect 48313 24850 48379 24853
rect 50200 24850 51000 24880
rect 48313 24848 51000 24850
rect 48313 24792 48318 24848
rect 48374 24792 51000 24848
rect 48313 24790 51000 24792
rect 48313 24787 48379 24790
rect 50200 24760 51000 24790
rect 15929 24714 15995 24717
rect 35985 24714 36051 24717
rect 15929 24712 36051 24714
rect 15929 24656 15934 24712
rect 15990 24656 35990 24712
rect 36046 24656 36051 24712
rect 15929 24654 36051 24656
rect 15929 24651 15995 24654
rect 35985 24651 36051 24654
rect 29085 24578 29151 24581
rect 28950 24576 29151 24578
rect 28950 24520 29090 24576
rect 29146 24520 29151 24576
rect 28950 24518 29151 24520
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 2773 24442 2839 24445
rect 28950 24442 29010 24518
rect 29085 24515 29151 24518
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 23430 24382 29010 24442
rect 11881 24306 11947 24309
rect 21081 24306 21147 24309
rect 11881 24304 21147 24306
rect 11881 24248 11886 24304
rect 11942 24248 21086 24304
rect 21142 24248 21147 24304
rect 11881 24246 21147 24248
rect 11881 24243 11947 24246
rect 21081 24243 21147 24246
rect 21357 24306 21423 24309
rect 23430 24306 23490 24382
rect 21357 24304 23490 24306
rect 21357 24248 21362 24304
rect 21418 24248 23490 24304
rect 21357 24246 23490 24248
rect 26141 24306 26207 24309
rect 29177 24306 29243 24309
rect 26141 24304 29243 24306
rect 26141 24248 26146 24304
rect 26202 24248 29182 24304
rect 29238 24248 29243 24304
rect 26141 24246 29243 24248
rect 21357 24243 21423 24246
rect 26141 24243 26207 24246
rect 29177 24243 29243 24246
rect 6545 24170 6611 24173
rect 24209 24170 24275 24173
rect 6545 24168 24275 24170
rect 6545 24112 6550 24168
rect 6606 24112 24214 24168
rect 24270 24112 24275 24168
rect 6545 24110 24275 24112
rect 6545 24107 6611 24110
rect 24209 24107 24275 24110
rect 24485 24170 24551 24173
rect 25313 24170 25379 24173
rect 24485 24168 25379 24170
rect 24485 24112 24490 24168
rect 24546 24112 25318 24168
rect 25374 24112 25379 24168
rect 24485 24110 25379 24112
rect 24485 24107 24551 24110
rect 25313 24107 25379 24110
rect 25497 24170 25563 24173
rect 41321 24170 41387 24173
rect 25497 24168 41387 24170
rect 25497 24112 25502 24168
rect 25558 24112 41326 24168
rect 41382 24112 41387 24168
rect 25497 24110 41387 24112
rect 25497 24107 25563 24110
rect 41321 24107 41387 24110
rect 0 24034 800 24064
rect 3509 24034 3575 24037
rect 0 24032 3575 24034
rect 0 23976 3514 24032
rect 3570 23976 3575 24032
rect 0 23974 3575 23976
rect 0 23944 800 23974
rect 3509 23971 3575 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 49509 23898 49575 23901
rect 50200 23898 51000 23928
rect 49509 23896 51000 23898
rect 49509 23840 49514 23896
rect 49570 23840 51000 23896
rect 49509 23838 51000 23840
rect 49509 23835 49575 23838
rect 50200 23808 51000 23838
rect 15101 23762 15167 23765
rect 17953 23762 18019 23765
rect 15101 23760 18019 23762
rect 15101 23704 15106 23760
rect 15162 23704 17958 23760
rect 18014 23704 18019 23760
rect 15101 23702 18019 23704
rect 15101 23699 15167 23702
rect 17953 23699 18019 23702
rect 18137 23762 18203 23765
rect 33869 23762 33935 23765
rect 18137 23760 33935 23762
rect 18137 23704 18142 23760
rect 18198 23704 33874 23760
rect 33930 23704 33935 23760
rect 18137 23702 33935 23704
rect 18137 23699 18203 23702
rect 33869 23699 33935 23702
rect 0 23626 800 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 800 23566
rect 4061 23563 4127 23566
rect 4654 23564 4660 23628
rect 4724 23626 4730 23628
rect 7189 23626 7255 23629
rect 4724 23624 7255 23626
rect 4724 23568 7194 23624
rect 7250 23568 7255 23624
rect 4724 23566 7255 23568
rect 4724 23564 4730 23566
rect 7189 23563 7255 23566
rect 12249 23626 12315 23629
rect 32121 23626 32187 23629
rect 12249 23624 32187 23626
rect 12249 23568 12254 23624
rect 12310 23568 32126 23624
rect 32182 23568 32187 23624
rect 12249 23566 32187 23568
rect 12249 23563 12315 23566
rect 32121 23563 32187 23566
rect 6729 23492 6795 23493
rect 6678 23490 6684 23492
rect 6638 23430 6684 23490
rect 6748 23488 6795 23492
rect 6790 23432 6795 23488
rect 6678 23428 6684 23430
rect 6748 23428 6795 23432
rect 6729 23427 6795 23428
rect 11881 23490 11947 23493
rect 22185 23492 22251 23493
rect 12014 23490 12020 23492
rect 11881 23488 12020 23490
rect 11881 23432 11886 23488
rect 11942 23432 12020 23488
rect 11881 23430 12020 23432
rect 11881 23427 11947 23430
rect 12014 23428 12020 23430
rect 12084 23428 12090 23492
rect 22134 23490 22140 23492
rect 22094 23430 22140 23490
rect 22204 23488 22251 23492
rect 22246 23432 22251 23488
rect 22134 23428 22140 23430
rect 22204 23428 22251 23432
rect 22185 23427 22251 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 0 23218 800 23248
rect 4061 23218 4127 23221
rect 0 23216 4127 23218
rect 0 23160 4066 23216
rect 4122 23160 4127 23216
rect 0 23158 4127 23160
rect 0 23128 800 23158
rect 4061 23155 4127 23158
rect 14457 23218 14523 23221
rect 24761 23218 24827 23221
rect 14457 23216 24827 23218
rect 14457 23160 14462 23216
rect 14518 23160 24766 23216
rect 24822 23160 24827 23216
rect 14457 23158 24827 23160
rect 14457 23155 14523 23158
rect 24761 23155 24827 23158
rect 14365 23082 14431 23085
rect 34513 23082 34579 23085
rect 14365 23080 34579 23082
rect 14365 23024 14370 23080
rect 14426 23024 34518 23080
rect 34574 23024 34579 23080
rect 14365 23022 34579 23024
rect 14365 23019 14431 23022
rect 34513 23019 34579 23022
rect 49325 22946 49391 22949
rect 50200 22946 51000 22976
rect 49325 22944 51000 22946
rect 49325 22888 49330 22944
rect 49386 22888 51000 22944
rect 49325 22886 51000 22888
rect 49325 22883 49391 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 50200 22856 51000 22886
rect 47946 22815 48262 22816
rect 3877 22810 3943 22813
rect 0 22808 3943 22810
rect 0 22752 3882 22808
rect 3938 22752 3943 22808
rect 0 22750 3943 22752
rect 0 22720 800 22750
rect 3877 22747 3943 22750
rect 11789 22810 11855 22813
rect 17401 22810 17467 22813
rect 27705 22810 27771 22813
rect 11789 22808 17467 22810
rect 11789 22752 11794 22808
rect 11850 22752 17406 22808
rect 17462 22752 17467 22808
rect 11789 22750 17467 22752
rect 11789 22747 11855 22750
rect 17401 22747 17467 22750
rect 18462 22808 27771 22810
rect 18462 22752 27710 22808
rect 27766 22752 27771 22808
rect 18462 22750 27771 22752
rect 15469 22674 15535 22677
rect 18462 22674 18522 22750
rect 27705 22747 27771 22750
rect 15469 22672 18522 22674
rect 15469 22616 15474 22672
rect 15530 22616 18522 22672
rect 15469 22614 18522 22616
rect 20621 22674 20687 22677
rect 32949 22674 33015 22677
rect 20621 22672 33015 22674
rect 20621 22616 20626 22672
rect 20682 22616 32954 22672
rect 33010 22616 33015 22672
rect 20621 22614 33015 22616
rect 15469 22611 15535 22614
rect 20621 22611 20687 22614
rect 32949 22611 33015 22614
rect 4153 22538 4219 22541
rect 17401 22538 17467 22541
rect 22553 22538 22619 22541
rect 24025 22538 24091 22541
rect 4153 22536 17234 22538
rect 4153 22480 4158 22536
rect 4214 22480 17234 22536
rect 4153 22478 17234 22480
rect 4153 22475 4219 22478
rect 0 22402 800 22432
rect 17174 22402 17234 22478
rect 17401 22536 22619 22538
rect 17401 22480 17406 22536
rect 17462 22480 22558 22536
rect 22614 22480 22619 22536
rect 17401 22478 22619 22480
rect 17401 22475 17467 22478
rect 22553 22475 22619 22478
rect 22694 22536 24091 22538
rect 22694 22480 24030 22536
rect 24086 22480 24091 22536
rect 22694 22478 24091 22480
rect 22694 22402 22754 22478
rect 24025 22475 24091 22478
rect 0 22342 2330 22402
rect 17174 22342 22754 22402
rect 0 22312 800 22342
rect 2270 22130 2330 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 17174 22206 22110 22266
rect 3509 22130 3575 22133
rect 2270 22128 3575 22130
rect 2270 22072 3514 22128
rect 3570 22072 3575 22128
rect 2270 22070 3575 22072
rect 3509 22067 3575 22070
rect 6637 22130 6703 22133
rect 17174 22130 17234 22206
rect 6637 22128 17234 22130
rect 6637 22072 6642 22128
rect 6698 22072 17234 22128
rect 6637 22070 17234 22072
rect 22050 22130 22110 22206
rect 23565 22130 23631 22133
rect 22050 22128 23631 22130
rect 22050 22072 23570 22128
rect 23626 22072 23631 22128
rect 22050 22070 23631 22072
rect 6637 22067 6703 22070
rect 23565 22067 23631 22070
rect 24393 22130 24459 22133
rect 26509 22130 26575 22133
rect 27429 22130 27495 22133
rect 24393 22128 27495 22130
rect 24393 22072 24398 22128
rect 24454 22072 26514 22128
rect 26570 22072 27434 22128
rect 27490 22072 27495 22128
rect 24393 22070 27495 22072
rect 24393 22067 24459 22070
rect 26509 22067 26575 22070
rect 27429 22067 27495 22070
rect 0 21994 800 22024
rect 3233 21994 3299 21997
rect 0 21992 3299 21994
rect 0 21936 3238 21992
rect 3294 21936 3299 21992
rect 0 21934 3299 21936
rect 0 21904 800 21934
rect 3233 21931 3299 21934
rect 16757 21994 16823 21997
rect 24577 21994 24643 21997
rect 39297 21994 39363 21997
rect 16757 21992 24643 21994
rect 16757 21936 16762 21992
rect 16818 21936 24582 21992
rect 24638 21936 24643 21992
rect 16757 21934 24643 21936
rect 16757 21931 16823 21934
rect 24577 21931 24643 21934
rect 26926 21992 39363 21994
rect 26926 21936 39302 21992
rect 39358 21936 39363 21992
rect 26926 21934 39363 21936
rect 20161 21858 20227 21861
rect 26926 21858 26986 21934
rect 39297 21931 39363 21934
rect 49509 21994 49575 21997
rect 50200 21994 51000 22024
rect 49509 21992 51000 21994
rect 49509 21936 49514 21992
rect 49570 21936 51000 21992
rect 49509 21934 51000 21936
rect 49509 21931 49575 21934
rect 50200 21904 51000 21934
rect 20161 21856 26986 21858
rect 20161 21800 20166 21856
rect 20222 21800 26986 21856
rect 20161 21798 26986 21800
rect 20161 21795 20227 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 18505 21722 18571 21725
rect 21265 21722 21331 21725
rect 18505 21720 21331 21722
rect 18505 21664 18510 21720
rect 18566 21664 21270 21720
rect 21326 21664 21331 21720
rect 18505 21662 21331 21664
rect 18505 21659 18571 21662
rect 21265 21659 21331 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 5625 21586 5691 21589
rect 6177 21586 6243 21589
rect 8661 21586 8727 21589
rect 5625 21584 8727 21586
rect 5625 21528 5630 21584
rect 5686 21528 6182 21584
rect 6238 21528 8666 21584
rect 8722 21528 8727 21584
rect 5625 21526 8727 21528
rect 5625 21523 5691 21526
rect 6177 21523 6243 21526
rect 8661 21523 8727 21526
rect 18413 21586 18479 21589
rect 30005 21586 30071 21589
rect 18413 21584 30071 21586
rect 18413 21528 18418 21584
rect 18474 21528 30010 21584
rect 30066 21528 30071 21584
rect 18413 21526 30071 21528
rect 18413 21523 18479 21526
rect 30005 21523 30071 21526
rect 10225 21450 10291 21453
rect 11237 21450 11303 21453
rect 15377 21450 15443 21453
rect 10225 21448 15443 21450
rect 10225 21392 10230 21448
rect 10286 21392 11242 21448
rect 11298 21392 15382 21448
rect 15438 21392 15443 21448
rect 10225 21390 15443 21392
rect 10225 21387 10291 21390
rect 11237 21387 11303 21390
rect 15377 21387 15443 21390
rect 15561 21450 15627 21453
rect 31109 21450 31175 21453
rect 15561 21448 31175 21450
rect 15561 21392 15566 21448
rect 15622 21392 31114 21448
rect 31170 21392 31175 21448
rect 15561 21390 31175 21392
rect 15561 21387 15627 21390
rect 31109 21387 31175 21390
rect 6862 21252 6868 21316
rect 6932 21314 6938 21316
rect 9765 21314 9831 21317
rect 6932 21312 9831 21314
rect 6932 21256 9770 21312
rect 9826 21256 9831 21312
rect 6932 21254 9831 21256
rect 6932 21252 6938 21254
rect 9765 21251 9831 21254
rect 17585 21314 17651 21317
rect 20345 21314 20411 21317
rect 17585 21312 20411 21314
rect 17585 21256 17590 21312
rect 17646 21256 20350 21312
rect 20406 21256 20411 21312
rect 17585 21254 20411 21256
rect 17585 21251 17651 21254
rect 20345 21251 20411 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 3969 21178 4035 21181
rect 11830 21178 11836 21180
rect 3969 21176 11836 21178
rect 3969 21120 3974 21176
rect 4030 21120 11836 21176
rect 3969 21118 11836 21120
rect 3969 21115 4035 21118
rect 11830 21116 11836 21118
rect 11900 21116 11906 21180
rect 13905 21178 13971 21181
rect 19057 21178 19123 21181
rect 13905 21176 19123 21178
rect 13905 21120 13910 21176
rect 13966 21120 19062 21176
rect 19118 21120 19123 21176
rect 13905 21118 19123 21120
rect 13905 21115 13971 21118
rect 19057 21115 19123 21118
rect 26417 21178 26483 21181
rect 27981 21178 28047 21181
rect 26417 21176 28047 21178
rect 26417 21120 26422 21176
rect 26478 21120 27986 21176
rect 28042 21120 28047 21176
rect 26417 21118 28047 21120
rect 26417 21115 26483 21118
rect 27981 21115 28047 21118
rect 4245 21042 4311 21045
rect 32029 21042 32095 21045
rect 4245 21040 32095 21042
rect 4245 20984 4250 21040
rect 4306 20984 32034 21040
rect 32090 20984 32095 21040
rect 4245 20982 32095 20984
rect 4245 20979 4311 20982
rect 32029 20979 32095 20982
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 8109 20906 8175 20909
rect 8518 20906 8524 20908
rect 8109 20904 8524 20906
rect 8109 20848 8114 20904
rect 8170 20848 8524 20904
rect 8109 20846 8524 20848
rect 8109 20843 8175 20846
rect 8518 20844 8524 20846
rect 8588 20844 8594 20908
rect 17401 20906 17467 20909
rect 28625 20906 28691 20909
rect 17401 20904 28691 20906
rect 17401 20848 17406 20904
rect 17462 20848 28630 20904
rect 28686 20848 28691 20904
rect 17401 20846 28691 20848
rect 17401 20843 17467 20846
rect 28625 20843 28691 20846
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 6126 20708 6132 20772
rect 6196 20770 6202 20772
rect 6269 20770 6335 20773
rect 6196 20768 6335 20770
rect 6196 20712 6274 20768
rect 6330 20712 6335 20768
rect 6196 20710 6335 20712
rect 6196 20708 6202 20710
rect 6269 20707 6335 20710
rect 11094 20708 11100 20772
rect 11164 20770 11170 20772
rect 11329 20770 11395 20773
rect 11164 20768 11395 20770
rect 11164 20712 11334 20768
rect 11390 20712 11395 20768
rect 11164 20710 11395 20712
rect 11164 20708 11170 20710
rect 11329 20707 11395 20710
rect 15745 20770 15811 20773
rect 17033 20772 17099 20773
rect 15878 20770 15884 20772
rect 15745 20768 15884 20770
rect 15745 20712 15750 20768
rect 15806 20712 15884 20768
rect 15745 20710 15884 20712
rect 15745 20707 15811 20710
rect 15878 20708 15884 20710
rect 15948 20708 15954 20772
rect 16982 20770 16988 20772
rect 16942 20710 16988 20770
rect 17052 20768 17099 20772
rect 17094 20712 17099 20768
rect 16982 20708 16988 20710
rect 17052 20708 17099 20712
rect 17033 20707 17099 20708
rect 22737 20770 22803 20773
rect 25681 20770 25747 20773
rect 22737 20768 25747 20770
rect 22737 20712 22742 20768
rect 22798 20712 25686 20768
rect 25742 20712 25747 20768
rect 22737 20710 25747 20712
rect 22737 20707 22803 20710
rect 25681 20707 25747 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 3601 20634 3667 20637
rect 7046 20634 7052 20636
rect 3601 20632 7052 20634
rect 3601 20576 3606 20632
rect 3662 20576 7052 20632
rect 3601 20574 7052 20576
rect 3601 20571 3667 20574
rect 7046 20572 7052 20574
rect 7116 20572 7122 20636
rect 18413 20634 18479 20637
rect 27521 20634 27587 20637
rect 18413 20632 27587 20634
rect 18413 20576 18418 20632
rect 18474 20576 27526 20632
rect 27582 20576 27587 20632
rect 18413 20574 27587 20576
rect 18413 20571 18479 20574
rect 27521 20571 27587 20574
rect 3601 20498 3667 20501
rect 9397 20498 9463 20501
rect 3601 20496 9463 20498
rect 3601 20440 3606 20496
rect 3662 20440 9402 20496
rect 9458 20440 9463 20496
rect 3601 20438 9463 20440
rect 3601 20435 3667 20438
rect 9397 20435 9463 20438
rect 16481 20498 16547 20501
rect 27705 20498 27771 20501
rect 46841 20498 46907 20501
rect 16481 20496 27771 20498
rect 16481 20440 16486 20496
rect 16542 20440 27710 20496
rect 27766 20440 27771 20496
rect 16481 20438 27771 20440
rect 16481 20435 16547 20438
rect 27705 20435 27771 20438
rect 31710 20496 46907 20498
rect 31710 20440 46846 20496
rect 46902 20440 46907 20496
rect 31710 20438 46907 20440
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 13629 20362 13695 20365
rect 13905 20362 13971 20365
rect 13629 20360 13971 20362
rect 13629 20304 13634 20360
rect 13690 20304 13910 20360
rect 13966 20304 13971 20360
rect 13629 20302 13971 20304
rect 13629 20299 13695 20302
rect 13905 20299 13971 20302
rect 17217 20362 17283 20365
rect 18413 20362 18479 20365
rect 30281 20362 30347 20365
rect 17217 20360 18479 20362
rect 17217 20304 17222 20360
rect 17278 20304 18418 20360
rect 18474 20304 18479 20360
rect 17217 20302 18479 20304
rect 17217 20299 17283 20302
rect 18413 20299 18479 20302
rect 22050 20360 30347 20362
rect 22050 20304 30286 20360
rect 30342 20304 30347 20360
rect 22050 20302 30347 20304
rect 13353 20226 13419 20229
rect 22050 20226 22110 20302
rect 30281 20299 30347 20302
rect 13353 20224 22110 20226
rect 13353 20168 13358 20224
rect 13414 20168 22110 20224
rect 13353 20166 22110 20168
rect 25313 20226 25379 20229
rect 31710 20226 31770 20438
rect 46841 20435 46907 20438
rect 25313 20224 31770 20226
rect 25313 20168 25318 20224
rect 25374 20168 31770 20224
rect 25313 20166 31770 20168
rect 13353 20163 13419 20166
rect 25313 20163 25379 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 13629 20090 13695 20093
rect 17125 20090 17191 20093
rect 13629 20088 17191 20090
rect 13629 20032 13634 20088
rect 13690 20032 17130 20088
rect 17186 20032 17191 20088
rect 13629 20030 17191 20032
rect 13629 20027 13695 20030
rect 17125 20027 17191 20030
rect 0 19954 800 19984
rect 1393 19954 1459 19957
rect 0 19952 1459 19954
rect 0 19896 1398 19952
rect 1454 19896 1459 19952
rect 0 19894 1459 19896
rect 0 19864 800 19894
rect 1393 19891 1459 19894
rect 5625 19954 5691 19957
rect 6545 19954 6611 19957
rect 28625 19954 28691 19957
rect 5625 19952 28691 19954
rect 5625 19896 5630 19952
rect 5686 19896 6550 19952
rect 6606 19896 28630 19952
rect 28686 19896 28691 19952
rect 5625 19894 28691 19896
rect 5625 19891 5691 19894
rect 6545 19891 6611 19894
rect 28625 19891 28691 19894
rect 11789 19818 11855 19821
rect 32397 19818 32463 19821
rect 11789 19816 32463 19818
rect 11789 19760 11794 19816
rect 11850 19760 32402 19816
rect 32458 19760 32463 19816
rect 11789 19758 32463 19760
rect 11789 19755 11855 19758
rect 32397 19755 32463 19758
rect 16798 19620 16804 19684
rect 16868 19682 16874 19684
rect 16941 19682 17007 19685
rect 17769 19682 17835 19685
rect 16868 19680 17835 19682
rect 16868 19624 16946 19680
rect 17002 19624 17774 19680
rect 17830 19624 17835 19680
rect 16868 19622 17835 19624
rect 16868 19620 16874 19622
rect 16941 19619 17007 19622
rect 17769 19619 17835 19622
rect 18505 19682 18571 19685
rect 25313 19682 25379 19685
rect 18505 19680 25379 19682
rect 18505 19624 18510 19680
rect 18566 19624 25318 19680
rect 25374 19624 25379 19680
rect 18505 19622 25379 19624
rect 18505 19619 18571 19622
rect 25313 19619 25379 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2957 19546 3023 19549
rect 0 19544 3023 19546
rect 0 19488 2962 19544
rect 3018 19488 3023 19544
rect 0 19486 3023 19488
rect 0 19456 800 19486
rect 2957 19483 3023 19486
rect 14365 19546 14431 19549
rect 15101 19546 15167 19549
rect 14365 19544 15167 19546
rect 14365 19488 14370 19544
rect 14426 19488 15106 19544
rect 15162 19488 15167 19544
rect 14365 19486 15167 19488
rect 14365 19483 14431 19486
rect 15101 19483 15167 19486
rect 20253 19546 20319 19549
rect 21633 19546 21699 19549
rect 27521 19546 27587 19549
rect 20253 19544 27587 19546
rect 20253 19488 20258 19544
rect 20314 19488 21638 19544
rect 21694 19488 27526 19544
rect 27582 19488 27587 19544
rect 20253 19486 27587 19488
rect 20253 19483 20319 19486
rect 21633 19483 21699 19486
rect 27521 19483 27587 19486
rect 5022 19348 5028 19412
rect 5092 19410 5098 19412
rect 5349 19410 5415 19413
rect 5092 19408 5415 19410
rect 5092 19352 5354 19408
rect 5410 19352 5415 19408
rect 5092 19350 5415 19352
rect 5092 19348 5098 19350
rect 5349 19347 5415 19350
rect 6453 19410 6519 19413
rect 7414 19410 7420 19412
rect 6453 19408 7420 19410
rect 6453 19352 6458 19408
rect 6514 19352 7420 19408
rect 6453 19350 7420 19352
rect 6453 19347 6519 19350
rect 7414 19348 7420 19350
rect 7484 19348 7490 19412
rect 10409 19410 10475 19413
rect 30649 19410 30715 19413
rect 10409 19408 30715 19410
rect 10409 19352 10414 19408
rect 10470 19352 30654 19408
rect 30710 19352 30715 19408
rect 10409 19350 30715 19352
rect 10409 19347 10475 19350
rect 30649 19347 30715 19350
rect 6913 19274 6979 19277
rect 19425 19274 19491 19277
rect 6913 19272 19491 19274
rect 6913 19216 6918 19272
rect 6974 19216 19430 19272
rect 19486 19216 19491 19272
rect 6913 19214 19491 19216
rect 6913 19211 6979 19214
rect 19425 19211 19491 19214
rect 25865 19274 25931 19277
rect 44449 19274 44515 19277
rect 25865 19272 44515 19274
rect 25865 19216 25870 19272
rect 25926 19216 44454 19272
rect 44510 19216 44515 19272
rect 25865 19214 44515 19216
rect 25865 19211 25931 19214
rect 44449 19211 44515 19214
rect 0 19138 800 19168
rect 2681 19138 2747 19141
rect 0 19136 2747 19138
rect 0 19080 2686 19136
rect 2742 19080 2747 19136
rect 0 19078 2747 19080
rect 0 19048 800 19078
rect 2681 19075 2747 19078
rect 17677 19138 17743 19141
rect 18229 19138 18295 19141
rect 17677 19136 18295 19138
rect 17677 19080 17682 19136
rect 17738 19080 18234 19136
rect 18290 19080 18295 19136
rect 17677 19078 18295 19080
rect 17677 19075 17743 19078
rect 18229 19075 18295 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 18638 19002 18644 19004
rect 14782 18942 18644 19002
rect 9765 18866 9831 18869
rect 14782 18866 14842 18942
rect 18638 18940 18644 18942
rect 18708 19002 18714 19004
rect 18708 18942 22110 19002
rect 18708 18940 18714 18942
rect 9765 18864 14842 18866
rect 9765 18808 9770 18864
rect 9826 18808 14842 18864
rect 9765 18806 14842 18808
rect 17125 18866 17191 18869
rect 18505 18866 18571 18869
rect 17125 18864 18571 18866
rect 17125 18808 17130 18864
rect 17186 18808 18510 18864
rect 18566 18808 18571 18864
rect 17125 18806 18571 18808
rect 22050 18866 22110 18942
rect 23841 18866 23907 18869
rect 43989 18866 44055 18869
rect 22050 18864 44055 18866
rect 22050 18808 23846 18864
rect 23902 18808 43994 18864
rect 44050 18808 44055 18864
rect 22050 18806 44055 18808
rect 9765 18803 9831 18806
rect 17125 18803 17191 18806
rect 18505 18803 18571 18806
rect 23841 18803 23907 18806
rect 43989 18803 44055 18806
rect 0 18730 800 18760
rect 2865 18730 2931 18733
rect 0 18728 2931 18730
rect 0 18672 2870 18728
rect 2926 18672 2931 18728
rect 0 18670 2931 18672
rect 0 18640 800 18670
rect 2865 18667 2931 18670
rect 10961 18730 11027 18733
rect 12341 18730 12407 18733
rect 10961 18728 12407 18730
rect 10961 18672 10966 18728
rect 11022 18672 12346 18728
rect 12402 18672 12407 18728
rect 10961 18670 12407 18672
rect 10961 18667 11027 18670
rect 12341 18667 12407 18670
rect 14181 18730 14247 18733
rect 16481 18730 16547 18733
rect 19701 18730 19767 18733
rect 35893 18730 35959 18733
rect 14181 18728 18476 18730
rect 14181 18672 14186 18728
rect 14242 18672 16486 18728
rect 16542 18672 18476 18728
rect 14181 18670 18476 18672
rect 14181 18667 14247 18670
rect 16481 18667 16547 18670
rect 10869 18594 10935 18597
rect 14733 18594 14799 18597
rect 10869 18592 14799 18594
rect 10869 18536 10874 18592
rect 10930 18536 14738 18592
rect 14794 18536 14799 18592
rect 10869 18534 14799 18536
rect 10869 18531 10935 18534
rect 14733 18531 14799 18534
rect 15009 18594 15075 18597
rect 15142 18594 15148 18596
rect 15009 18592 15148 18594
rect 15009 18536 15014 18592
rect 15070 18536 15148 18592
rect 15009 18534 15148 18536
rect 15009 18531 15075 18534
rect 15142 18532 15148 18534
rect 15212 18532 15218 18596
rect 18416 18594 18476 18670
rect 19701 18728 35959 18730
rect 19701 18672 19706 18728
rect 19762 18672 35898 18728
rect 35954 18672 35959 18728
rect 19701 18670 35959 18672
rect 19701 18667 19767 18670
rect 35893 18667 35959 18670
rect 19977 18594 20043 18597
rect 18416 18592 20043 18594
rect 18416 18536 19982 18592
rect 20038 18536 20043 18592
rect 18416 18534 20043 18536
rect 19977 18531 20043 18534
rect 22829 18594 22895 18597
rect 26693 18594 26759 18597
rect 22829 18592 26759 18594
rect 22829 18536 22834 18592
rect 22890 18536 26698 18592
rect 26754 18536 26759 18592
rect 22829 18534 26759 18536
rect 22829 18531 22895 18534
rect 26693 18531 26759 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 9489 18458 9555 18461
rect 11881 18458 11947 18461
rect 9489 18456 11947 18458
rect 9489 18400 9494 18456
rect 9550 18400 11886 18456
rect 11942 18400 11947 18456
rect 9489 18398 11947 18400
rect 9489 18395 9555 18398
rect 11881 18395 11947 18398
rect 18689 18458 18755 18461
rect 26141 18458 26207 18461
rect 18689 18456 26207 18458
rect 18689 18400 18694 18456
rect 18750 18400 26146 18456
rect 26202 18400 26207 18456
rect 18689 18398 26207 18400
rect 18689 18395 18755 18398
rect 26141 18395 26207 18398
rect 0 18322 800 18352
rect 2773 18322 2839 18325
rect 12433 18322 12499 18325
rect 0 18320 2839 18322
rect 0 18264 2778 18320
rect 2834 18264 2839 18320
rect 0 18262 2839 18264
rect 0 18232 800 18262
rect 2773 18259 2839 18262
rect 7606 18320 12499 18322
rect 7606 18264 12438 18320
rect 12494 18264 12499 18320
rect 7606 18262 12499 18264
rect 2681 18186 2747 18189
rect 7606 18186 7666 18262
rect 12433 18259 12499 18262
rect 15101 18322 15167 18325
rect 27613 18322 27679 18325
rect 15101 18320 27679 18322
rect 15101 18264 15106 18320
rect 15162 18264 27618 18320
rect 27674 18264 27679 18320
rect 15101 18262 27679 18264
rect 15101 18259 15167 18262
rect 27613 18259 27679 18262
rect 2681 18184 7666 18186
rect 2681 18128 2686 18184
rect 2742 18128 7666 18184
rect 2681 18126 7666 18128
rect 12157 18186 12223 18189
rect 31661 18186 31727 18189
rect 12157 18184 31727 18186
rect 12157 18128 12162 18184
rect 12218 18128 31666 18184
rect 31722 18128 31727 18184
rect 12157 18126 31727 18128
rect 2681 18123 2747 18126
rect 12157 18123 12223 18126
rect 31661 18123 31727 18126
rect 7189 18050 7255 18053
rect 9213 18050 9279 18053
rect 7189 18048 9279 18050
rect 7189 17992 7194 18048
rect 7250 17992 9218 18048
rect 9274 17992 9279 18048
rect 7189 17990 9279 17992
rect 7189 17987 7255 17990
rect 9213 17987 9279 17990
rect 14549 18050 14615 18053
rect 18689 18050 18755 18053
rect 14549 18048 18755 18050
rect 14549 17992 14554 18048
rect 14610 17992 18694 18048
rect 18750 17992 18755 18048
rect 14549 17990 18755 17992
rect 14549 17987 14615 17990
rect 18689 17987 18755 17990
rect 19425 18050 19491 18053
rect 21909 18050 21975 18053
rect 19425 18048 21975 18050
rect 19425 17992 19430 18048
rect 19486 17992 21914 18048
rect 21970 17992 21975 18048
rect 19425 17990 21975 17992
rect 19425 17987 19491 17990
rect 21909 17987 21975 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 3601 17914 3667 17917
rect 5625 17914 5691 17917
rect 3601 17912 5691 17914
rect 3601 17856 3606 17912
rect 3662 17856 5630 17912
rect 5686 17856 5691 17912
rect 3601 17854 5691 17856
rect 3601 17851 3667 17854
rect 5625 17851 5691 17854
rect 6269 17914 6335 17917
rect 9581 17914 9647 17917
rect 6269 17912 9647 17914
rect 6269 17856 6274 17912
rect 6330 17856 9586 17912
rect 9642 17856 9647 17912
rect 6269 17854 9647 17856
rect 6269 17851 6335 17854
rect 9581 17851 9647 17854
rect 13537 17914 13603 17917
rect 20069 17914 20135 17917
rect 13537 17912 20135 17914
rect 13537 17856 13542 17912
rect 13598 17856 20074 17912
rect 20130 17856 20135 17912
rect 13537 17854 20135 17856
rect 13537 17851 13603 17854
rect 20069 17851 20135 17854
rect 27521 17914 27587 17917
rect 30649 17914 30715 17917
rect 27521 17912 30715 17914
rect 27521 17856 27526 17912
rect 27582 17856 30654 17912
rect 30710 17856 30715 17912
rect 27521 17854 30715 17856
rect 27521 17851 27587 17854
rect 30649 17851 30715 17854
rect 4429 17778 4495 17781
rect 14457 17778 14523 17781
rect 4429 17776 14523 17778
rect 4429 17720 4434 17776
rect 4490 17720 14462 17776
rect 14518 17720 14523 17776
rect 4429 17718 14523 17720
rect 4429 17715 4495 17718
rect 14457 17715 14523 17718
rect 19977 17778 20043 17781
rect 24209 17778 24275 17781
rect 30189 17778 30255 17781
rect 19977 17776 30255 17778
rect 19977 17720 19982 17776
rect 20038 17720 24214 17776
rect 24270 17720 30194 17776
rect 30250 17720 30255 17776
rect 19977 17718 30255 17720
rect 19977 17715 20043 17718
rect 24209 17715 24275 17718
rect 30189 17715 30255 17718
rect 6545 17642 6611 17645
rect 12065 17642 12131 17645
rect 6545 17640 12131 17642
rect 6545 17584 6550 17640
rect 6606 17584 12070 17640
rect 12126 17584 12131 17640
rect 6545 17582 12131 17584
rect 6545 17579 6611 17582
rect 12065 17579 12131 17582
rect 14089 17642 14155 17645
rect 20161 17642 20227 17645
rect 14089 17640 20227 17642
rect 14089 17584 14094 17640
rect 14150 17584 20166 17640
rect 20222 17584 20227 17640
rect 14089 17582 20227 17584
rect 14089 17579 14155 17582
rect 20161 17579 20227 17582
rect 24393 17642 24459 17645
rect 30097 17642 30163 17645
rect 24393 17640 30163 17642
rect 24393 17584 24398 17640
rect 24454 17584 30102 17640
rect 30158 17584 30163 17640
rect 24393 17582 30163 17584
rect 24393 17579 24459 17582
rect 30097 17579 30163 17582
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 1761 17370 1827 17373
rect 6453 17370 6519 17373
rect 1761 17368 6519 17370
rect 1761 17312 1766 17368
rect 1822 17312 6458 17368
rect 6514 17312 6519 17368
rect 1761 17310 6519 17312
rect 1761 17307 1827 17310
rect 6453 17307 6519 17310
rect 9949 17370 10015 17373
rect 12893 17370 12959 17373
rect 9949 17368 12959 17370
rect 9949 17312 9954 17368
rect 10010 17312 12898 17368
rect 12954 17312 12959 17368
rect 9949 17310 12959 17312
rect 9949 17307 10015 17310
rect 12893 17307 12959 17310
rect 18781 17370 18847 17373
rect 18965 17370 19031 17373
rect 23565 17370 23631 17373
rect 18781 17368 23631 17370
rect 18781 17312 18786 17368
rect 18842 17312 18970 17368
rect 19026 17312 23570 17368
rect 23626 17312 23631 17368
rect 18781 17310 23631 17312
rect 18781 17307 18847 17310
rect 18965 17307 19031 17310
rect 23565 17307 23631 17310
rect 5349 17234 5415 17237
rect 9765 17234 9831 17237
rect 5349 17232 9831 17234
rect 5349 17176 5354 17232
rect 5410 17176 9770 17232
rect 9826 17176 9831 17232
rect 5349 17174 9831 17176
rect 5349 17171 5415 17174
rect 9765 17171 9831 17174
rect 11053 17234 11119 17237
rect 19241 17234 19307 17237
rect 11053 17232 19307 17234
rect 11053 17176 11058 17232
rect 11114 17176 19246 17232
rect 19302 17176 19307 17232
rect 11053 17174 19307 17176
rect 11053 17171 11119 17174
rect 19241 17171 19307 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 5901 17098 5967 17101
rect 6545 17098 6611 17101
rect 5901 17096 6611 17098
rect 5901 17040 5906 17096
rect 5962 17040 6550 17096
rect 6606 17040 6611 17096
rect 5901 17038 6611 17040
rect 5901 17035 5967 17038
rect 6545 17035 6611 17038
rect 9029 17098 9095 17101
rect 26601 17098 26667 17101
rect 9029 17096 26667 17098
rect 9029 17040 9034 17096
rect 9090 17040 26606 17096
rect 26662 17040 26667 17096
rect 9029 17038 26667 17040
rect 9029 17035 9095 17038
rect 26601 17035 26667 17038
rect 7046 16900 7052 16964
rect 7116 16962 7122 16964
rect 11145 16962 11211 16965
rect 7116 16960 11211 16962
rect 7116 16904 11150 16960
rect 11206 16904 11211 16960
rect 7116 16902 11211 16904
rect 7116 16900 7122 16902
rect 11145 16899 11211 16902
rect 13813 16962 13879 16965
rect 18454 16962 18460 16964
rect 13813 16960 18460 16962
rect 13813 16904 13818 16960
rect 13874 16904 18460 16960
rect 13813 16902 18460 16904
rect 13813 16899 13879 16902
rect 18454 16900 18460 16902
rect 18524 16900 18530 16964
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 4705 16826 4771 16829
rect 8017 16826 8083 16829
rect 4705 16824 8083 16826
rect 4705 16768 4710 16824
rect 4766 16768 8022 16824
rect 8078 16768 8083 16824
rect 4705 16766 8083 16768
rect 4705 16763 4771 16766
rect 8017 16763 8083 16766
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 2865 16690 2931 16693
rect 5441 16690 5507 16693
rect 2865 16688 5507 16690
rect 2865 16632 2870 16688
rect 2926 16632 5446 16688
rect 5502 16632 5507 16688
rect 2865 16630 5507 16632
rect 2865 16627 2931 16630
rect 5441 16627 5507 16630
rect 6453 16690 6519 16693
rect 8109 16690 8175 16693
rect 6453 16688 8175 16690
rect 6453 16632 6458 16688
rect 6514 16632 8114 16688
rect 8170 16632 8175 16688
rect 6453 16630 8175 16632
rect 6453 16627 6519 16630
rect 8109 16627 8175 16630
rect 12433 16690 12499 16693
rect 29545 16690 29611 16693
rect 12433 16688 29611 16690
rect 12433 16632 12438 16688
rect 12494 16632 29550 16688
rect 29606 16632 29611 16688
rect 12433 16630 29611 16632
rect 12433 16627 12499 16630
rect 29545 16627 29611 16630
rect 4521 16554 4587 16557
rect 6085 16554 6151 16557
rect 6729 16554 6795 16557
rect 4521 16552 6795 16554
rect 4521 16496 4526 16552
rect 4582 16496 6090 16552
rect 6146 16496 6734 16552
rect 6790 16496 6795 16552
rect 4521 16494 6795 16496
rect 4521 16491 4587 16494
rect 6085 16491 6151 16494
rect 6729 16491 6795 16494
rect 7465 16554 7531 16557
rect 11053 16554 11119 16557
rect 7465 16552 11119 16554
rect 7465 16496 7470 16552
rect 7526 16496 11058 16552
rect 11114 16496 11119 16552
rect 7465 16494 11119 16496
rect 7465 16491 7531 16494
rect 11053 16491 11119 16494
rect 14365 16554 14431 16557
rect 28533 16554 28599 16557
rect 14365 16552 28599 16554
rect 14365 16496 14370 16552
rect 14426 16496 28538 16552
rect 28594 16496 28599 16552
rect 14365 16494 28599 16496
rect 14365 16491 14431 16494
rect 28533 16491 28599 16494
rect 12198 16356 12204 16420
rect 12268 16418 12274 16420
rect 13629 16418 13695 16421
rect 12268 16416 13695 16418
rect 12268 16360 13634 16416
rect 13690 16360 13695 16416
rect 12268 16358 13695 16360
rect 12268 16356 12274 16358
rect 13629 16355 13695 16358
rect 15142 16356 15148 16420
rect 15212 16418 15218 16420
rect 15377 16418 15443 16421
rect 15212 16416 15443 16418
rect 15212 16360 15382 16416
rect 15438 16360 15443 16416
rect 15212 16358 15443 16360
rect 15212 16356 15218 16358
rect 15377 16355 15443 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 12065 16282 12131 16285
rect 17125 16282 17191 16285
rect 12065 16280 17191 16282
rect 12065 16224 12070 16280
rect 12126 16224 17130 16280
rect 17186 16224 17191 16280
rect 12065 16222 17191 16224
rect 12065 16219 12131 16222
rect 17125 16219 17191 16222
rect 18454 16220 18460 16284
rect 18524 16282 18530 16284
rect 22921 16282 22987 16285
rect 18524 16280 22987 16282
rect 18524 16224 22926 16280
rect 22982 16224 22987 16280
rect 18524 16222 22987 16224
rect 18524 16220 18530 16222
rect 22921 16219 22987 16222
rect 2037 16146 2103 16149
rect 8385 16146 8451 16149
rect 2037 16144 8451 16146
rect 2037 16088 2042 16144
rect 2098 16088 8390 16144
rect 8446 16088 8451 16144
rect 2037 16086 8451 16088
rect 2037 16083 2103 16086
rect 8385 16083 8451 16086
rect 10041 16146 10107 16149
rect 10317 16146 10383 16149
rect 10041 16144 10383 16146
rect 10041 16088 10046 16144
rect 10102 16088 10322 16144
rect 10378 16088 10383 16144
rect 10041 16086 10383 16088
rect 10041 16083 10107 16086
rect 10317 16083 10383 16086
rect 10869 16146 10935 16149
rect 21265 16146 21331 16149
rect 10869 16144 21331 16146
rect 10869 16088 10874 16144
rect 10930 16088 21270 16144
rect 21326 16088 21331 16144
rect 10869 16086 21331 16088
rect 10869 16083 10935 16086
rect 21265 16083 21331 16086
rect 21817 16146 21883 16149
rect 25129 16146 25195 16149
rect 21817 16144 25195 16146
rect 21817 16088 21822 16144
rect 21878 16088 25134 16144
rect 25190 16088 25195 16144
rect 21817 16086 25195 16088
rect 21817 16083 21883 16086
rect 25129 16083 25195 16086
rect 8477 16010 8543 16013
rect 9857 16010 9923 16013
rect 8477 16008 9923 16010
rect 8477 15952 8482 16008
rect 8538 15952 9862 16008
rect 9918 15952 9923 16008
rect 8477 15950 9923 15952
rect 8477 15947 8543 15950
rect 9857 15947 9923 15950
rect 10961 16010 11027 16013
rect 28993 16010 29059 16013
rect 10961 16008 29059 16010
rect 10961 15952 10966 16008
rect 11022 15952 28998 16008
rect 29054 15952 29059 16008
rect 10961 15950 29059 15952
rect 10961 15947 11027 15950
rect 28993 15947 29059 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 5717 15874 5783 15877
rect 6545 15874 6611 15877
rect 9673 15874 9739 15877
rect 5717 15872 9739 15874
rect 5717 15816 5722 15872
rect 5778 15816 6550 15872
rect 6606 15816 9678 15872
rect 9734 15816 9739 15872
rect 5717 15814 9739 15816
rect 5717 15811 5783 15814
rect 6545 15811 6611 15814
rect 9673 15811 9739 15814
rect 16941 15874 17007 15877
rect 20253 15874 20319 15877
rect 16941 15872 20319 15874
rect 16941 15816 16946 15872
rect 17002 15816 20258 15872
rect 20314 15816 20319 15872
rect 16941 15814 20319 15816
rect 16941 15811 17007 15814
rect 20253 15811 20319 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 7557 15738 7623 15741
rect 9489 15738 9555 15741
rect 7557 15736 9555 15738
rect 7557 15680 7562 15736
rect 7618 15680 9494 15736
rect 9550 15680 9555 15736
rect 7557 15678 9555 15680
rect 7557 15675 7623 15678
rect 9489 15675 9555 15678
rect 13353 15738 13419 15741
rect 19701 15738 19767 15741
rect 13353 15736 19767 15738
rect 13353 15680 13358 15736
rect 13414 15680 19706 15736
rect 19762 15680 19767 15736
rect 13353 15678 19767 15680
rect 13353 15675 13419 15678
rect 19701 15675 19767 15678
rect 6637 15602 6703 15605
rect 8661 15602 8727 15605
rect 6637 15600 8727 15602
rect 6637 15544 6642 15600
rect 6698 15544 8666 15600
rect 8722 15544 8727 15600
rect 6637 15542 8727 15544
rect 6637 15539 6703 15542
rect 8661 15539 8727 15542
rect 9213 15600 9279 15605
rect 9213 15544 9218 15600
rect 9274 15544 9279 15600
rect 9213 15539 9279 15544
rect 12065 15602 12131 15605
rect 29913 15602 29979 15605
rect 12065 15600 29979 15602
rect 12065 15544 12070 15600
rect 12126 15544 29918 15600
rect 29974 15544 29979 15600
rect 12065 15542 29979 15544
rect 12065 15539 12131 15542
rect 29913 15539 29979 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 7189 15466 7255 15469
rect 9216 15466 9276 15539
rect 7189 15464 9276 15466
rect 7189 15408 7194 15464
rect 7250 15408 9276 15464
rect 7189 15406 9276 15408
rect 9857 15466 9923 15469
rect 31937 15466 32003 15469
rect 9857 15464 32003 15466
rect 9857 15408 9862 15464
rect 9918 15408 31942 15464
rect 31998 15408 32003 15464
rect 9857 15406 32003 15408
rect 7189 15403 7255 15406
rect 9857 15403 9923 15406
rect 31937 15403 32003 15406
rect 1393 15330 1459 15333
rect 7649 15330 7715 15333
rect 1393 15328 7715 15330
rect 1393 15272 1398 15328
rect 1454 15272 7654 15328
rect 7710 15272 7715 15328
rect 1393 15270 7715 15272
rect 1393 15267 1459 15270
rect 7649 15267 7715 15270
rect 11053 15330 11119 15333
rect 16021 15330 16087 15333
rect 11053 15328 16087 15330
rect 11053 15272 11058 15328
rect 11114 15272 16026 15328
rect 16082 15272 16087 15328
rect 11053 15270 16087 15272
rect 11053 15267 11119 15270
rect 16021 15267 16087 15270
rect 20529 15330 20595 15333
rect 25589 15330 25655 15333
rect 20529 15328 25655 15330
rect 20529 15272 20534 15328
rect 20590 15272 25594 15328
rect 25650 15272 25655 15328
rect 20529 15270 25655 15272
rect 20529 15267 20595 15270
rect 25589 15267 25655 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 9857 15194 9923 15197
rect 10961 15194 11027 15197
rect 13077 15194 13143 15197
rect 9857 15192 13143 15194
rect 9857 15136 9862 15192
rect 9918 15136 10966 15192
rect 11022 15136 13082 15192
rect 13138 15136 13143 15192
rect 9857 15134 13143 15136
rect 9857 15131 9923 15134
rect 10961 15131 11027 15134
rect 13077 15131 13143 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 4061 15058 4127 15061
rect 4429 15058 4495 15061
rect 4061 15056 4495 15058
rect 4061 15000 4066 15056
rect 4122 15000 4434 15056
rect 4490 15000 4495 15056
rect 4061 14998 4495 15000
rect 4061 14995 4127 14998
rect 4429 14995 4495 14998
rect 6177 15058 6243 15061
rect 7833 15058 7899 15061
rect 11973 15058 12039 15061
rect 33409 15058 33475 15061
rect 6177 15056 10978 15058
rect 6177 15000 6182 15056
rect 6238 15000 7838 15056
rect 7894 15000 10978 15056
rect 6177 14998 10978 15000
rect 6177 14995 6243 14998
rect 7833 14995 7899 14998
rect 3509 14922 3575 14925
rect 7649 14922 7715 14925
rect 3509 14920 7715 14922
rect 3509 14864 3514 14920
rect 3570 14864 7654 14920
rect 7710 14864 7715 14920
rect 3509 14862 7715 14864
rect 10918 14922 10978 14998
rect 11973 15056 33475 15058
rect 11973 15000 11978 15056
rect 12034 15000 33414 15056
rect 33470 15000 33475 15056
rect 11973 14998 33475 15000
rect 11973 14995 12039 14998
rect 33409 14995 33475 14998
rect 11329 14922 11395 14925
rect 10918 14920 11395 14922
rect 10918 14864 11334 14920
rect 11390 14864 11395 14920
rect 10918 14862 11395 14864
rect 3509 14859 3575 14862
rect 7649 14859 7715 14862
rect 11329 14859 11395 14862
rect 14733 14922 14799 14925
rect 15837 14922 15903 14925
rect 14733 14920 15903 14922
rect 14733 14864 14738 14920
rect 14794 14864 15842 14920
rect 15898 14864 15903 14920
rect 14733 14862 15903 14864
rect 14733 14859 14799 14862
rect 15837 14859 15903 14862
rect 17125 14922 17191 14925
rect 19333 14922 19399 14925
rect 17125 14920 19399 14922
rect 17125 14864 17130 14920
rect 17186 14864 19338 14920
rect 19394 14864 19399 14920
rect 17125 14862 19399 14864
rect 17125 14859 17191 14862
rect 19333 14859 19399 14862
rect 5533 14786 5599 14789
rect 8753 14786 8819 14789
rect 5533 14784 8819 14786
rect 5533 14728 5538 14784
rect 5594 14728 8758 14784
rect 8814 14728 8819 14784
rect 5533 14726 8819 14728
rect 5533 14723 5599 14726
rect 8753 14723 8819 14726
rect 10041 14786 10107 14789
rect 12065 14786 12131 14789
rect 10041 14784 12131 14786
rect 10041 14728 10046 14784
rect 10102 14728 12070 14784
rect 12126 14728 12131 14784
rect 10041 14726 12131 14728
rect 10041 14723 10107 14726
rect 12065 14723 12131 14726
rect 15561 14786 15627 14789
rect 18781 14786 18847 14789
rect 15561 14784 18847 14786
rect 15561 14728 15566 14784
rect 15622 14728 18786 14784
rect 18842 14728 18847 14784
rect 15561 14726 18847 14728
rect 15561 14723 15627 14726
rect 18781 14723 18847 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 5165 14650 5231 14653
rect 8569 14650 8635 14653
rect 5165 14648 8635 14650
rect 5165 14592 5170 14648
rect 5226 14592 8574 14648
rect 8630 14592 8635 14648
rect 5165 14590 8635 14592
rect 5165 14587 5231 14590
rect 8569 14587 8635 14590
rect 5717 14514 5783 14517
rect 9489 14514 9555 14517
rect 5717 14512 9555 14514
rect 5717 14456 5722 14512
rect 5778 14456 9494 14512
rect 9550 14456 9555 14512
rect 5717 14454 9555 14456
rect 5717 14451 5783 14454
rect 9489 14451 9555 14454
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 2589 14106 2655 14109
rect 3550 14106 3556 14108
rect 2589 14104 3556 14106
rect 2589 14048 2594 14104
rect 2650 14048 3556 14104
rect 2589 14046 3556 14048
rect 2589 14043 2655 14046
rect 3550 14044 3556 14046
rect 3620 14044 3626 14108
rect 1761 13970 1827 13973
rect 20069 13970 20135 13973
rect 1761 13968 20135 13970
rect 1761 13912 1766 13968
rect 1822 13912 20074 13968
rect 20130 13912 20135 13968
rect 1761 13910 20135 13912
rect 1761 13907 1827 13910
rect 20069 13907 20135 13910
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 10777 13834 10843 13837
rect 13905 13834 13971 13837
rect 10777 13832 13971 13834
rect 10777 13776 10782 13832
rect 10838 13776 13910 13832
rect 13966 13776 13971 13832
rect 10777 13774 13971 13776
rect 10777 13771 10843 13774
rect 13905 13771 13971 13774
rect 4705 13698 4771 13701
rect 6862 13698 6868 13700
rect 4705 13696 6868 13698
rect 4705 13640 4710 13696
rect 4766 13640 6868 13696
rect 4705 13638 6868 13640
rect 4705 13635 4771 13638
rect 6862 13636 6868 13638
rect 6932 13636 6938 13700
rect 7230 13636 7236 13700
rect 7300 13698 7306 13700
rect 11094 13698 11100 13700
rect 7300 13638 11100 13698
rect 7300 13636 7306 13638
rect 11094 13636 11100 13638
rect 11164 13636 11170 13700
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 4245 13562 4311 13565
rect 9489 13562 9555 13565
rect 4245 13560 9555 13562
rect 4245 13504 4250 13560
rect 4306 13504 9494 13560
rect 9550 13504 9555 13560
rect 4245 13502 9555 13504
rect 4245 13499 4311 13502
rect 9489 13499 9555 13502
rect 17125 13562 17191 13565
rect 17493 13562 17559 13565
rect 18505 13562 18571 13565
rect 17125 13560 18571 13562
rect 17125 13504 17130 13560
rect 17186 13504 17498 13560
rect 17554 13504 18510 13560
rect 18566 13504 18571 13560
rect 17125 13502 18571 13504
rect 17125 13499 17191 13502
rect 17493 13499 17559 13502
rect 18505 13499 18571 13502
rect 0 13426 800 13456
rect 1301 13426 1367 13429
rect 0 13424 1367 13426
rect 0 13368 1306 13424
rect 1362 13368 1367 13424
rect 0 13366 1367 13368
rect 0 13336 800 13366
rect 1301 13363 1367 13366
rect 9397 13426 9463 13429
rect 31017 13426 31083 13429
rect 9397 13424 31083 13426
rect 9397 13368 9402 13424
rect 9458 13368 31022 13424
rect 31078 13368 31083 13424
rect 9397 13366 31083 13368
rect 9397 13363 9463 13366
rect 31017 13363 31083 13366
rect 3325 13290 3391 13293
rect 22277 13290 22343 13293
rect 3325 13288 22343 13290
rect 3325 13232 3330 13288
rect 3386 13232 22282 13288
rect 22338 13232 22343 13288
rect 3325 13230 22343 13232
rect 3325 13227 3391 13230
rect 22277 13227 22343 13230
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 3601 13018 3667 13021
rect 0 13016 3667 13018
rect 0 12960 3606 13016
rect 3662 12960 3667 13016
rect 0 12958 3667 12960
rect 0 12928 800 12958
rect 3601 12955 3667 12958
rect 11605 13018 11671 13021
rect 17769 13018 17835 13021
rect 11605 13016 17835 13018
rect 11605 12960 11610 13016
rect 11666 12960 17774 13016
rect 17830 12960 17835 13016
rect 11605 12958 17835 12960
rect 11605 12955 11671 12958
rect 17769 12955 17835 12958
rect 7097 12884 7163 12885
rect 7046 12820 7052 12884
rect 7116 12882 7163 12884
rect 10685 12882 10751 12885
rect 22093 12882 22159 12885
rect 7116 12880 7208 12882
rect 7158 12824 7208 12880
rect 7116 12822 7208 12824
rect 10685 12880 22159 12882
rect 10685 12824 10690 12880
rect 10746 12824 22098 12880
rect 22154 12824 22159 12880
rect 10685 12822 22159 12824
rect 7116 12820 7163 12822
rect 7097 12819 7163 12820
rect 10685 12819 10751 12822
rect 22093 12819 22159 12822
rect 12985 12746 13051 12749
rect 17769 12746 17835 12749
rect 20897 12746 20963 12749
rect 26141 12746 26207 12749
rect 12985 12744 17602 12746
rect 12985 12688 12990 12744
rect 13046 12688 17602 12744
rect 12985 12686 17602 12688
rect 12985 12683 13051 12686
rect 0 12610 800 12640
rect 1669 12610 1735 12613
rect 0 12608 1735 12610
rect 0 12552 1674 12608
rect 1730 12552 1735 12608
rect 0 12550 1735 12552
rect 0 12520 800 12550
rect 1669 12547 1735 12550
rect 7189 12610 7255 12613
rect 7741 12610 7807 12613
rect 7189 12608 7807 12610
rect 7189 12552 7194 12608
rect 7250 12552 7746 12608
rect 7802 12552 7807 12608
rect 7189 12550 7807 12552
rect 17542 12610 17602 12686
rect 17769 12744 26207 12746
rect 17769 12688 17774 12744
rect 17830 12688 20902 12744
rect 20958 12688 26146 12744
rect 26202 12688 26207 12744
rect 17769 12686 26207 12688
rect 17769 12683 17835 12686
rect 20897 12683 20963 12686
rect 26141 12683 26207 12686
rect 17769 12610 17835 12613
rect 17542 12608 17835 12610
rect 17542 12552 17774 12608
rect 17830 12552 17835 12608
rect 17542 12550 17835 12552
rect 7189 12547 7255 12550
rect 7741 12547 7807 12550
rect 17769 12547 17835 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 4153 12474 4219 12477
rect 12014 12474 12020 12476
rect 4153 12472 12020 12474
rect 4153 12416 4158 12472
rect 4214 12416 12020 12472
rect 4153 12414 12020 12416
rect 4153 12411 4219 12414
rect 12014 12412 12020 12414
rect 12084 12412 12090 12476
rect 12525 12338 12591 12341
rect 19149 12338 19215 12341
rect 12525 12336 19215 12338
rect 12525 12280 12530 12336
rect 12586 12280 19154 12336
rect 19210 12280 19215 12336
rect 12525 12278 19215 12280
rect 12525 12275 12591 12278
rect 19149 12275 19215 12278
rect 0 12202 800 12232
rect 1301 12202 1367 12205
rect 0 12200 1367 12202
rect 0 12144 1306 12200
rect 1362 12144 1367 12200
rect 0 12142 1367 12144
rect 0 12112 800 12142
rect 1301 12139 1367 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 14181 11930 14247 11933
rect 15193 11930 15259 11933
rect 18597 11932 18663 11933
rect 18597 11930 18644 11932
rect 14181 11928 15259 11930
rect 14181 11872 14186 11928
rect 14242 11872 15198 11928
rect 15254 11872 15259 11928
rect 14181 11870 15259 11872
rect 18552 11928 18644 11930
rect 18552 11872 18602 11928
rect 18552 11870 18644 11872
rect 14181 11867 14247 11870
rect 15193 11867 15259 11870
rect 18597 11868 18644 11870
rect 18708 11868 18714 11932
rect 18597 11867 18663 11868
rect 0 11794 800 11824
rect 1577 11794 1643 11797
rect 0 11792 1643 11794
rect 0 11736 1582 11792
rect 1638 11736 1643 11792
rect 0 11734 1643 11736
rect 0 11704 800 11734
rect 1577 11731 1643 11734
rect 8201 11794 8267 11797
rect 8753 11794 8819 11797
rect 8201 11792 8819 11794
rect 8201 11736 8206 11792
rect 8262 11736 8758 11792
rect 8814 11736 8819 11792
rect 8201 11734 8819 11736
rect 8201 11731 8267 11734
rect 8753 11731 8819 11734
rect 11830 11732 11836 11796
rect 11900 11794 11906 11796
rect 11973 11794 12039 11797
rect 11900 11792 12039 11794
rect 11900 11736 11978 11792
rect 12034 11736 12039 11792
rect 11900 11734 12039 11736
rect 11900 11732 11906 11734
rect 11973 11731 12039 11734
rect 9765 11658 9831 11661
rect 13445 11658 13511 11661
rect 9765 11656 13511 11658
rect 9765 11600 9770 11656
rect 9826 11600 13450 11656
rect 13506 11600 13511 11656
rect 9765 11598 13511 11600
rect 9765 11595 9831 11598
rect 13445 11595 13511 11598
rect 4981 11524 5047 11525
rect 4981 11520 5028 11524
rect 5092 11522 5098 11524
rect 7005 11522 7071 11525
rect 7414 11522 7420 11524
rect 4981 11464 4986 11520
rect 4981 11460 5028 11464
rect 5092 11462 5138 11522
rect 7005 11520 7420 11522
rect 7005 11464 7010 11520
rect 7066 11464 7420 11520
rect 7005 11462 7420 11464
rect 5092 11460 5098 11462
rect 4981 11459 5047 11460
rect 7005 11459 7071 11462
rect 7414 11460 7420 11462
rect 7484 11460 7490 11524
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 4889 11386 4955 11389
rect 9765 11386 9831 11389
rect 0 11326 2790 11386
rect 0 11296 800 11326
rect 2730 11250 2790 11326
rect 4889 11384 9831 11386
rect 4889 11328 4894 11384
rect 4950 11328 9770 11384
rect 9826 11328 9831 11384
rect 4889 11326 9831 11328
rect 4889 11323 4955 11326
rect 9765 11323 9831 11326
rect 3325 11250 3391 11253
rect 2730 11248 3391 11250
rect 2730 11192 3330 11248
rect 3386 11192 3391 11248
rect 2730 11190 3391 11192
rect 3325 11187 3391 11190
rect 3601 11250 3667 11253
rect 11053 11250 11119 11253
rect 16798 11250 16804 11252
rect 3601 11248 9506 11250
rect 3601 11192 3606 11248
rect 3662 11192 9506 11248
rect 3601 11190 9506 11192
rect 3601 11187 3667 11190
rect 6177 11116 6243 11117
rect 6126 11114 6132 11116
rect 6086 11054 6132 11114
rect 6196 11112 6243 11116
rect 6238 11056 6243 11112
rect 6126 11052 6132 11054
rect 6196 11052 6243 11056
rect 8518 11052 8524 11116
rect 8588 11114 8594 11116
rect 9305 11114 9371 11117
rect 8588 11112 9371 11114
rect 8588 11056 9310 11112
rect 9366 11056 9371 11112
rect 8588 11054 9371 11056
rect 9446 11114 9506 11190
rect 11053 11248 16804 11250
rect 11053 11192 11058 11248
rect 11114 11192 16804 11248
rect 11053 11190 16804 11192
rect 11053 11187 11119 11190
rect 16798 11188 16804 11190
rect 16868 11188 16874 11252
rect 28901 11114 28967 11117
rect 9446 11112 28967 11114
rect 9446 11056 28906 11112
rect 28962 11056 28967 11112
rect 9446 11054 28967 11056
rect 8588 11052 8594 11054
rect 6177 11051 6243 11052
rect 9305 11051 9371 11054
rect 28901 11051 28967 11054
rect 0 10978 800 11008
rect 2773 10978 2839 10981
rect 0 10976 2839 10978
rect 0 10920 2778 10976
rect 2834 10920 2839 10976
rect 0 10918 2839 10920
rect 0 10888 800 10918
rect 2773 10915 2839 10918
rect 10225 10978 10291 10981
rect 12198 10978 12204 10980
rect 10225 10976 12204 10978
rect 10225 10920 10230 10976
rect 10286 10920 12204 10976
rect 10225 10918 12204 10920
rect 10225 10915 10291 10918
rect 12198 10916 12204 10918
rect 12268 10916 12274 10980
rect 17309 10978 17375 10981
rect 17769 10978 17835 10981
rect 17309 10976 17835 10978
rect 17309 10920 17314 10976
rect 17370 10920 17774 10976
rect 17830 10920 17835 10976
rect 17309 10918 17835 10920
rect 17309 10915 17375 10918
rect 17769 10915 17835 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 7281 10706 7347 10709
rect 16982 10706 16988 10708
rect 7281 10704 16988 10706
rect 7281 10648 7286 10704
rect 7342 10648 16988 10704
rect 7281 10646 16988 10648
rect 7281 10643 7347 10646
rect 16982 10644 16988 10646
rect 17052 10644 17058 10708
rect 0 10570 800 10600
rect 3601 10570 3667 10573
rect 0 10568 3667 10570
rect 0 10512 3606 10568
rect 3662 10512 3667 10568
rect 0 10510 3667 10512
rect 0 10480 800 10510
rect 3601 10507 3667 10510
rect 5349 10570 5415 10573
rect 22134 10570 22140 10572
rect 5349 10568 22140 10570
rect 5349 10512 5354 10568
rect 5410 10512 22140 10568
rect 5349 10510 22140 10512
rect 5349 10507 5415 10510
rect 22134 10508 22140 10510
rect 22204 10508 22210 10572
rect 6361 10434 6427 10437
rect 6678 10434 6684 10436
rect 6361 10432 6684 10434
rect 6361 10376 6366 10432
rect 6422 10376 6684 10432
rect 6361 10374 6684 10376
rect 6361 10371 6427 10374
rect 6678 10372 6684 10374
rect 6748 10372 6754 10436
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 2865 10162 2931 10165
rect 0 10160 2931 10162
rect 0 10104 2870 10160
rect 2926 10104 2931 10160
rect 0 10102 2931 10104
rect 0 10072 800 10102
rect 2865 10099 2931 10102
rect 4061 10026 4127 10029
rect 15878 10026 15884 10028
rect 4061 10024 15884 10026
rect 4061 9968 4066 10024
rect 4122 9968 15884 10024
rect 4061 9966 15884 9968
rect 4061 9963 4127 9966
rect 15878 9964 15884 9966
rect 15948 9964 15954 10028
rect 15285 9890 15351 9893
rect 16481 9890 16547 9893
rect 15285 9888 16547 9890
rect 15285 9832 15290 9888
rect 15346 9832 16486 9888
rect 16542 9832 16547 9888
rect 15285 9830 16547 9832
rect 15285 9827 15351 9830
rect 16481 9827 16547 9830
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 3601 9620 3667 9621
rect 3550 9556 3556 9620
rect 3620 9618 3667 9620
rect 4521 9618 4587 9621
rect 4654 9618 4660 9620
rect 3620 9616 3712 9618
rect 3662 9560 3712 9616
rect 3620 9558 3712 9560
rect 4521 9616 4660 9618
rect 4521 9560 4526 9616
rect 4582 9560 4660 9616
rect 4521 9558 4660 9560
rect 3620 9556 3667 9558
rect 3601 9555 3667 9556
rect 4521 9555 4587 9558
rect 4654 9556 4660 9558
rect 4724 9556 4730 9620
rect 0 9346 800 9376
rect 2497 9346 2563 9349
rect 0 9344 2563 9346
rect 0 9288 2502 9344
rect 2558 9288 2563 9344
rect 0 9286 2563 9288
rect 0 9256 800 9286
rect 2497 9283 2563 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 7189 9212 7255 9213
rect 7189 9210 7236 9212
rect 7144 9208 7236 9210
rect 7144 9152 7194 9208
rect 7144 9150 7236 9152
rect 7189 9148 7236 9150
rect 7300 9148 7306 9212
rect 7189 9147 7255 9148
rect 7741 9074 7807 9077
rect 23657 9074 23723 9077
rect 7741 9072 23723 9074
rect 7741 9016 7746 9072
rect 7802 9016 23662 9072
rect 23718 9016 23723 9072
rect 7741 9014 23723 9016
rect 7741 9011 7807 9014
rect 23657 9011 23723 9014
rect 0 8938 800 8968
rect 1761 8938 1827 8941
rect 0 8936 1827 8938
rect 0 8880 1766 8936
rect 1822 8880 1827 8936
rect 0 8878 1827 8880
rect 0 8848 800 8878
rect 1761 8875 1827 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 2865 8530 2931 8533
rect 0 8528 2931 8530
rect 0 8472 2870 8528
rect 2926 8472 2931 8528
rect 0 8470 2931 8472
rect 0 8440 800 8470
rect 2865 8467 2931 8470
rect 9581 8394 9647 8397
rect 32765 8394 32831 8397
rect 9581 8392 32831 8394
rect 9581 8336 9586 8392
rect 9642 8336 32770 8392
rect 32826 8336 32831 8392
rect 9581 8334 32831 8336
rect 9581 8331 9647 8334
rect 32765 8331 32831 8334
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 2405 8122 2471 8125
rect 0 8120 2471 8122
rect 0 8064 2410 8120
rect 2466 8064 2471 8120
rect 0 8062 2471 8064
rect 0 8032 800 8062
rect 2405 8059 2471 8062
rect 0 7714 800 7744
rect 3693 7714 3759 7717
rect 0 7712 3759 7714
rect 0 7656 3698 7712
rect 3754 7656 3759 7712
rect 0 7654 3759 7656
rect 0 7624 800 7654
rect 3693 7651 3759 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 0 7306 800 7336
rect 2865 7306 2931 7309
rect 0 7304 2931 7306
rect 0 7248 2870 7304
rect 2926 7248 2931 7304
rect 0 7246 2931 7248
rect 0 7216 800 7246
rect 2865 7243 2931 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 0 4450 800 4480
rect 1761 4450 1827 4453
rect 3509 4450 3575 4453
rect 0 4448 3575 4450
rect 0 4392 1766 4448
rect 1822 4392 3514 4448
rect 3570 4392 3575 4448
rect 0 4390 3575 4392
rect 0 4360 800 4390
rect 1761 4387 1827 4390
rect 3509 4387 3575 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 2681 4178 2747 4181
rect 6269 4178 6335 4181
rect 2681 4176 6335 4178
rect 2681 4120 2686 4176
rect 2742 4120 6274 4176
rect 6330 4120 6335 4176
rect 2681 4118 6335 4120
rect 2681 4115 2747 4118
rect 6269 4115 6335 4118
rect 0 4042 800 4072
rect 2865 4042 2931 4045
rect 0 4040 2931 4042
rect 0 3984 2870 4040
rect 2926 3984 2931 4040
rect 0 3982 2931 3984
rect 0 3952 800 3982
rect 2865 3979 2931 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 2773 2002 2839 2005
rect 0 2000 2839 2002
rect 0 1944 2778 2000
rect 2834 1944 2839 2000
rect 0 1942 2839 1944
rect 0 1912 800 1942
rect 2773 1939 2839 1942
rect 0 1594 800 1624
rect 3325 1594 3391 1597
rect 0 1592 3391 1594
rect 0 1536 3330 1592
rect 3386 1536 3391 1592
rect 0 1534 3391 1536
rect 0 1504 800 1534
rect 3325 1531 3391 1534
<< via3 >>
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 4660 23564 4724 23628
rect 6684 23488 6748 23492
rect 6684 23432 6734 23488
rect 6734 23432 6748 23488
rect 6684 23428 6748 23432
rect 12020 23428 12084 23492
rect 22140 23488 22204 23492
rect 22140 23432 22190 23488
rect 22190 23432 22204 23488
rect 22140 23428 22204 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 6868 21252 6932 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 11836 21116 11900 21180
rect 8524 20844 8588 20908
rect 6132 20708 6196 20772
rect 11100 20708 11164 20772
rect 15884 20708 15948 20772
rect 16988 20768 17052 20772
rect 16988 20712 17038 20768
rect 17038 20712 17052 20768
rect 16988 20708 17052 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 7052 20572 7116 20636
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 16804 19620 16868 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 5028 19348 5092 19412
rect 7420 19348 7484 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 18644 18940 18708 19004
rect 15148 18532 15212 18596
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 7052 16900 7116 16964
rect 18460 16900 18524 16964
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 12204 16356 12268 16420
rect 15148 16356 15212 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 18460 16220 18524 16284
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 3556 14044 3620 14108
rect 6868 13636 6932 13700
rect 7236 13636 7300 13700
rect 11100 13636 11164 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 7052 12880 7116 12884
rect 7052 12824 7102 12880
rect 7102 12824 7116 12880
rect 7052 12820 7116 12824
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 12020 12412 12084 12476
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 18644 11928 18708 11932
rect 18644 11872 18658 11928
rect 18658 11872 18708 11928
rect 18644 11868 18708 11872
rect 11836 11732 11900 11796
rect 5028 11520 5092 11524
rect 5028 11464 5042 11520
rect 5042 11464 5092 11520
rect 5028 11460 5092 11464
rect 7420 11460 7484 11524
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 6132 11112 6196 11116
rect 6132 11056 6182 11112
rect 6182 11056 6196 11112
rect 6132 11052 6196 11056
rect 8524 11052 8588 11116
rect 16804 11188 16868 11252
rect 12204 10916 12268 10980
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 16988 10644 17052 10708
rect 22140 10508 22204 10572
rect 6684 10372 6748 10436
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 15884 9964 15948 10028
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 3556 9616 3620 9620
rect 3556 9560 3606 9616
rect 3606 9560 3620 9616
rect 3556 9556 3620 9560
rect 4660 9556 4724 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7236 9208 7300 9212
rect 7236 9152 7250 9208
rect 7250 9152 7300 9208
rect 7236 9148 7300 9152
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 4659 23628 4725 23629
rect 4659 23564 4660 23628
rect 4724 23564 4725 23628
rect 4659 23563 4725 23564
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 3555 14108 3621 14109
rect 3555 14044 3556 14108
rect 3620 14044 3621 14108
rect 3555 14043 3621 14044
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 3558 9621 3618 14043
rect 4662 9621 4722 23563
rect 6683 23492 6749 23493
rect 6683 23428 6684 23492
rect 6748 23428 6749 23492
rect 6683 23427 6749 23428
rect 6131 20772 6197 20773
rect 6131 20708 6132 20772
rect 6196 20708 6197 20772
rect 6131 20707 6197 20708
rect 5027 19412 5093 19413
rect 5027 19348 5028 19412
rect 5092 19348 5093 19412
rect 5027 19347 5093 19348
rect 5030 11525 5090 19347
rect 5027 11524 5093 11525
rect 5027 11460 5028 11524
rect 5092 11460 5093 11524
rect 5027 11459 5093 11460
rect 6134 11117 6194 20707
rect 6131 11116 6197 11117
rect 6131 11052 6132 11116
rect 6196 11052 6197 11116
rect 6131 11051 6197 11052
rect 6686 10437 6746 23427
rect 7944 22880 8264 23904
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12019 23492 12085 23493
rect 12019 23428 12020 23492
rect 12084 23428 12085 23492
rect 12019 23427 12085 23428
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 6867 21316 6933 21317
rect 6867 21252 6868 21316
rect 6932 21252 6933 21316
rect 6867 21251 6933 21252
rect 6870 13701 6930 21251
rect 7944 20704 8264 21728
rect 11835 21180 11901 21181
rect 11835 21116 11836 21180
rect 11900 21116 11901 21180
rect 11835 21115 11901 21116
rect 8523 20908 8589 20909
rect 8523 20844 8524 20908
rect 8588 20844 8589 20908
rect 8523 20843 8589 20844
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7051 20636 7117 20637
rect 7051 20572 7052 20636
rect 7116 20572 7117 20636
rect 7051 20571 7117 20572
rect 7054 16965 7114 20571
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7419 19412 7485 19413
rect 7419 19348 7420 19412
rect 7484 19348 7485 19412
rect 7419 19347 7485 19348
rect 7051 16964 7117 16965
rect 7051 16900 7052 16964
rect 7116 16900 7117 16964
rect 7051 16899 7117 16900
rect 6867 13700 6933 13701
rect 6867 13636 6868 13700
rect 6932 13636 6933 13700
rect 6867 13635 6933 13636
rect 7054 12885 7114 16899
rect 7235 13700 7301 13701
rect 7235 13636 7236 13700
rect 7300 13636 7301 13700
rect 7235 13635 7301 13636
rect 7051 12884 7117 12885
rect 7051 12820 7052 12884
rect 7116 12820 7117 12884
rect 7051 12819 7117 12820
rect 6683 10436 6749 10437
rect 6683 10372 6684 10436
rect 6748 10372 6749 10436
rect 6683 10371 6749 10372
rect 3555 9620 3621 9621
rect 3555 9556 3556 9620
rect 3620 9556 3621 9620
rect 3555 9555 3621 9556
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 7238 9213 7298 13635
rect 7422 11525 7482 19347
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7419 11524 7485 11525
rect 7419 11460 7420 11524
rect 7484 11460 7485 11524
rect 7419 11459 7485 11460
rect 7944 10912 8264 11936
rect 8526 11117 8586 20843
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 11102 13701 11162 20707
rect 11099 13700 11165 13701
rect 11099 13636 11100 13700
rect 11164 13636 11165 13700
rect 11099 13635 11165 13636
rect 11838 11797 11898 21115
rect 12022 12477 12082 23427
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22139 23492 22205 23493
rect 22139 23428 22140 23492
rect 22204 23428 22205 23492
rect 22139 23427 22205 23428
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 16987 20772 17053 20773
rect 16987 20708 16988 20772
rect 17052 20708 17053 20772
rect 16987 20707 17053 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 15147 18596 15213 18597
rect 15147 18532 15148 18596
rect 15212 18532 15213 18596
rect 15147 18531 15213 18532
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12203 16420 12269 16421
rect 12203 16356 12204 16420
rect 12268 16356 12269 16420
rect 12203 16355 12269 16356
rect 12019 12476 12085 12477
rect 12019 12412 12020 12476
rect 12084 12412 12085 12476
rect 12019 12411 12085 12412
rect 11835 11796 11901 11797
rect 11835 11732 11836 11796
rect 11900 11732 11901 11796
rect 11835 11731 11901 11732
rect 8523 11116 8589 11117
rect 8523 11052 8524 11116
rect 8588 11052 8589 11116
rect 8523 11051 8589 11052
rect 12206 10981 12266 16355
rect 12944 15808 13264 16832
rect 15150 16421 15210 18531
rect 15147 16420 15213 16421
rect 15147 16356 15148 16420
rect 15212 16356 15213 16420
rect 15147 16355 15213 16356
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12203 10980 12269 10981
rect 12203 10916 12204 10980
rect 12268 10916 12269 10980
rect 12203 10915 12269 10916
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7235 9212 7301 9213
rect 7235 9148 7236 9212
rect 7300 9148 7301 9212
rect 7235 9147 7301 9148
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 15886 10029 15946 20707
rect 16803 19684 16869 19685
rect 16803 19620 16804 19684
rect 16868 19620 16869 19684
rect 16803 19619 16869 19620
rect 16806 11253 16866 19619
rect 16803 11252 16869 11253
rect 16803 11188 16804 11252
rect 16868 11188 16869 11252
rect 16803 11187 16869 11188
rect 16990 10709 17050 20707
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 18643 19004 18709 19005
rect 18643 18940 18644 19004
rect 18708 18940 18709 19004
rect 18643 18939 18709 18940
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 18459 16964 18525 16965
rect 18459 16900 18460 16964
rect 18524 16900 18525 16964
rect 18459 16899 18525 16900
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 18462 16285 18522 16899
rect 18459 16284 18525 16285
rect 18459 16220 18460 16284
rect 18524 16220 18525 16284
rect 18459 16219 18525 16220
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 18646 11933 18706 18939
rect 18643 11932 18709 11933
rect 18643 11868 18644 11932
rect 18708 11868 18709 11932
rect 18643 11867 18709 11868
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 16987 10708 17053 10709
rect 16987 10644 16988 10708
rect 17052 10644 17053 10708
rect 16987 10643 17053 10644
rect 15883 10028 15949 10029
rect 15883 9964 15884 10028
rect 15948 9964 15949 10028
rect 15883 9963 15949 9964
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 9824 18264 10848
rect 22142 10573 22202 23427
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22139 10572 22205 10573
rect 22139 10508 22140 10572
rect 22204 10508 22205 10572
rect 22139 10507 22205 10508
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1676037725
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 10672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 3404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 6072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 4232 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1676037725
transform 1 0 2208 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _134_
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _135_
timestamp 1676037725
transform 1 0 3404 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 33764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 32292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 33028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _147_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _149_
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1676037725
transform 1 0 18584 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _151_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1676037725
transform 1 0 33580 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1676037725
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 12328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 10120 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 10672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 35972 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 6624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 13616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 13800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 15364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1676037725
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1676037725
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1676037725
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1676037725
transform 1 0 3404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1676037725
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1676037725
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1676037725
transform 1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 32108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 31832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 34868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 3220 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 13064 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1676037725
transform 1 0 28336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 11132 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 4140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 34684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 32752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 33396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 35328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 33672 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 36616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 33028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 36984 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 37904 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 36800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 37260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 38180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 38916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 39836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 41768 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 41768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 31740 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 30912 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 30820 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 31924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 49036 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 43148 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 44804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 49220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14996 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30728 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27600 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 31464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 30912 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 30544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5336 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5428 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9568 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4232 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 6808 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10856 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28612 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 26956 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25760 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22172 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 14720 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 13616 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19596 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 24932 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1676037725
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1676037725
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1676037725
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1676037725
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_395
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_407
timestamp 1676037725
transform 1 0 38548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_22
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_28
timestamp 1676037725
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_40
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1676037725
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_142
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1676037725
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp 1676037725
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1676037725
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_116
timestamp 1676037725
transform 1 0 11776 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_28
timestamp 1676037725
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1676037725
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1676037725
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1676037725
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_205
timestamp 1676037725
transform 1 0 19964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_217
timestamp 1676037725
transform 1 0 21068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_229
timestamp 1676037725
transform 1 0 22172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1676037725
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1676037725
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1676037725
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1676037725
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1676037725
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_238
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1676037725
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1676037725
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1676037725
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_199
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_211
timestamp 1676037725
transform 1 0 20516 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1676037725
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1676037725
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1676037725
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1676037725
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_234
timestamp 1676037725
transform 1 0 22632 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_246
timestamp 1676037725
transform 1 0 23736 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_258
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_270
timestamp 1676037725
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1676037725
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1676037725
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1676037725
transform 1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_33
timestamp 1676037725
transform 1 0 4140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_45
timestamp 1676037725
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_57
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_69
timestamp 1676037725
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1676037725
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_106
timestamp 1676037725
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1676037725
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1676037725
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1676037725
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_127
timestamp 1676037725
transform 1 0 12788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_8
timestamp 1676037725
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1676037725
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_31
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_36
timestamp 1676037725
transform 1 0 4416 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_48
timestamp 1676037725
transform 1 0 5520 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_60
timestamp 1676037725
transform 1 0 6624 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_72
timestamp 1676037725
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1676037725
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_101
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_107
timestamp 1676037725
transform 1 0 10948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_128
timestamp 1676037725
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_169
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_181
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1676037725
transform 1 0 3128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1676037725
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_45
timestamp 1676037725
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_73
timestamp 1676037725
transform 1 0 7820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1676037725
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1676037725
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1676037725
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_129
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1676037725
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1676037725
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_34
timestamp 1676037725
transform 1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_42
timestamp 1676037725
transform 1 0 4968 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1676037725
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1676037725
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1676037725
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1676037725
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1676037725
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1676037725
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_19
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1676037725
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1676037725
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1676037725
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1676037725
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1676037725
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_294
timestamp 1676037725
transform 1 0 28152 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_298
timestamp 1676037725
transform 1 0 28520 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_310
timestamp 1676037725
transform 1 0 29624 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_322
timestamp 1676037725
transform 1 0 30728 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1676037725
transform 1 0 4048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_50
timestamp 1676037725
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1676037725
transform 1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1676037725
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1676037725
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1676037725
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1676037725
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_223
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_235
timestamp 1676037725
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_43
timestamp 1676037725
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1676037725
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1676037725
transform 1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1676037725
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_229
timestamp 1676037725
transform 1 0 22172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1676037725
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_265
timestamp 1676037725
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1676037725
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 1676037725
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1676037725
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1676037725
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1676037725
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1676037725
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1676037725
transform 1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1676037725
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1676037725
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1676037725
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1676037725
transform 1 0 31832 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_5
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_21
timestamp 1676037725
transform 1 0 3036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1676037725
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1676037725
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1676037725
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1676037725
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1676037725
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1676037725
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_228
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1676037725
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_255
timestamp 1676037725
transform 1 0 24564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1676037725
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_34
timestamp 1676037725
transform 1 0 4232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_42
timestamp 1676037725
transform 1 0 4968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_143
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1676037725
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_191
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1676037725
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_255
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_267
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_279
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 1676037725
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1676037725
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1676037725
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1676037725
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_19
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1676037725
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1676037725
transform 1 0 4508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_61
timestamp 1676037725
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1676037725
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1676037725
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_174
timestamp 1676037725
transform 1 0 17112 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1676037725
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_231
timestamp 1676037725
transform 1 0 22356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1676037725
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1676037725
transform 1 0 6348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_201
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_266
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1676037725
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1676037725
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1676037725
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1676037725
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_171
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_227
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1676037725
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1676037725
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1676037725
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1676037725
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1676037725
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_87
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_220
timestamp 1676037725
transform 1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1676037725
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1676037725
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_283
timestamp 1676037725
transform 1 0 27140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_295
timestamp 1676037725
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1676037725
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1676037725
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1676037725
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1676037725
transform 1 0 3404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1676037725
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1676037725
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1676037725
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_171
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_211
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1676037725
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_257
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_283
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_295
timestamp 1676037725
transform 1 0 28244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_307
timestamp 1676037725
transform 1 0 29348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1676037725
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1676037725
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1676037725
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1676037725
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_132
timestamp 1676037725
transform 1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1676037725
transform 1 0 19688 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_232
timestamp 1676037725
transform 1 0 22448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_237
timestamp 1676037725
transform 1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_255
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1676037725
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1676037725
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1676037725
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1676037725
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_173
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1676037725
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1676037725
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1676037725
transform 1 0 24104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_256
timestamp 1676037725
transform 1 0 24656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_283
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1676037725
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_290
timestamp 1676037725
transform 1 0 27784 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_302
timestamp 1676037725
transform 1 0 28888 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_314
timestamp 1676037725
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1676037725
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1676037725
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_123
timestamp 1676037725
transform 1 0 12420 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_160
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1676037725
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1676037725
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1676037725
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1676037725
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_88
timestamp 1676037725
transform 1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1676037725
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1676037725
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_150
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1676037725
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1676037725
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 1676037725
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_250
timestamp 1676037725
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_276
timestamp 1676037725
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1676037725
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_314
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_326
timestamp 1676037725
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_25
timestamp 1676037725
transform 1 0 3404 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1676037725
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1676037725
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1676037725
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1676037725
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_255
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1676037725
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1676037725
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1676037725
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1676037725
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1676037725
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 1676037725
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1676037725
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1676037725
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1676037725
transform 1 0 12788 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1676037725
transform 1 0 13156 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1676037725
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_230
timestamp 1676037725
transform 1 0 22264 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1676037725
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1676037725
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_286
timestamp 1676037725
transform 1 0 27416 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1676037725
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_25
timestamp 1676037725
transform 1 0 3404 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1676037725
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_99
timestamp 1676037725
transform 1 0 10212 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_103
timestamp 1676037725
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1676037725
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_216
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1676037725
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_324
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_336
timestamp 1676037725
transform 1 0 32016 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_348
timestamp 1676037725
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1676037725
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1676037725
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_135
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1676037725
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1676037725
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_274
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1676037725
transform 1 0 27416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_290
timestamp 1676037725
transform 1 0 27784 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_315
timestamp 1676037725
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_322
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1676037725
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1676037725
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_166
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1676037725
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1676037725
transform 1 0 23184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_293
timestamp 1676037725
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_314
timestamp 1676037725
transform 1 0 29992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_331
timestamp 1676037725
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_343
timestamp 1676037725
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1676037725
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1676037725
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_80
timestamp 1676037725
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_182
timestamp 1676037725
transform 1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_250
timestamp 1676037725
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_276
timestamp 1676037725
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1676037725
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1676037725
transform 1 0 5244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_108
timestamp 1676037725
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_114
timestamp 1676037725
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_144
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1676037725
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_226
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_269
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1676037725
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_344
timestamp 1676037725
transform 1 0 32752 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_356
timestamp 1676037725
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_61
timestamp 1676037725
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_67
timestamp 1676037725
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_91
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_129
timestamp 1676037725
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1676037725
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_330
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_343
timestamp 1676037725
transform 1 0 32660 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_355
timestamp 1676037725
transform 1 0 33764 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_367
timestamp 1676037725
transform 1 0 34868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_379
timestamp 1676037725
transform 1 0 35972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_507
timestamp 1676037725
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_25
timestamp 1676037725
transform 1 0 3404 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_57
timestamp 1676037725
transform 1 0 6348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1676037725
transform 1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_100
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1676037725
transform 1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1676037725
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_231
timestamp 1676037725
transform 1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1676037725
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_302
timestamp 1676037725
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_313
timestamp 1676037725
transform 1 0 29900 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_336
timestamp 1676037725
transform 1 0 32016 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_339
timestamp 1676037725
transform 1 0 32292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_352
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1676037725
transform 1 0 14260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_230
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1676037725
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1676037725
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1676037725
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1676037725
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_343
timestamp 1676037725
transform 1 0 32660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_351
timestamp 1676037725
transform 1 0 33396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_363
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_369
timestamp 1676037725
transform 1 0 35052 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1676037725
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_419
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_423
timestamp 1676037725
transform 1 0 40020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_435
timestamp 1676037725
transform 1 0 41124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_519
timestamp 1676037725
transform 1 0 48852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_25
timestamp 1676037725
transform 1 0 3404 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_87
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1676037725
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1676037725
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_281
timestamp 1676037725
transform 1 0 26956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_304
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_331
timestamp 1676037725
transform 1 0 31556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_337
timestamp 1676037725
transform 1 0 32108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_343
timestamp 1676037725
transform 1 0 32660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_351
timestamp 1676037725
transform 1 0 33396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_359
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_370
timestamp 1676037725
transform 1 0 35144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_384
timestamp 1676037725
transform 1 0 36432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_390
timestamp 1676037725
transform 1 0 36984 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_395
timestamp 1676037725
transform 1 0 37444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_407
timestamp 1676037725
transform 1 0 38548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1676037725
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1676037725
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1676037725
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_318
timestamp 1676037725
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_326
timestamp 1676037725
transform 1 0 31096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_331
timestamp 1676037725
transform 1 0 31556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_342
timestamp 1676037725
transform 1 0 32568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_353
timestamp 1676037725
transform 1 0 33580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_360
timestamp 1676037725
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_368
timestamp 1676037725
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_376
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_383
timestamp 1676037725
transform 1 0 36340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_395
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_401
timestamp 1676037725
transform 1 0 37996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_407
timestamp 1676037725
transform 1 0 38548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_413
timestamp 1676037725
transform 1 0 39100 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_423
timestamp 1676037725
transform 1 0 40020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_435
timestamp 1676037725
transform 1 0 41124 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_459
timestamp 1676037725
transform 1 0 43332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_465
timestamp 1676037725
transform 1 0 43884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_477
timestamp 1676037725
transform 1 0 44988 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_487
timestamp 1676037725
transform 1 0 45908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_495
timestamp 1676037725
transform 1 0 46644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_507
timestamp 1676037725
transform 1 0 47748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_511
timestamp 1676037725
transform 1 0 48116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_299
timestamp 1676037725
transform 1 0 28612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_325
timestamp 1676037725
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_331
timestamp 1676037725
transform 1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_346
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1676037725
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_371
timestamp 1676037725
transform 1 0 35236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_379
timestamp 1676037725
transform 1 0 35972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_386
timestamp 1676037725
transform 1 0 36616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_398
timestamp 1676037725
transform 1 0 37720 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_402
timestamp 1676037725
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_409
timestamp 1676037725
transform 1 0 38732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1676037725
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_440
timestamp 1676037725
transform 1 0 41584 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_444
timestamp 1676037725
transform 1 0 41952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_471
timestamp 1676037725
transform 1 0 44436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_519
timestamp 1676037725
transform 1 0 48852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_523
timestamp 1676037725
transform 1 0 49220 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 48392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 35512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 36064 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 37720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 41308 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 41308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 28336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1676037725
transform 1 0 42596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 44252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 49036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 48300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18676 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27232 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4600 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__194
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11224 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18492 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__195
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__196
timestamp 1676037725
transform 1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__197
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28336 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__198
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30084 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__188
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__189
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__169
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__175
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__176
timestamp 1676037725
transform 1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__177
timestamp 1676037725
transform 1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__178
timestamp 1676037725
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 30452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4140 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 32936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32568 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__187
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset_top_in
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable_top_in
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 17526 6188 17526 6188 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 15686 6222 15686 6222 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 14812 5746 14812 5746 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 13662 9639 13662 9639 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20838 17714 20838 17714 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 9752 10166 9752 10166 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 12558 13872 12558 13872 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 10580 13838 10580 13838 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 8602 9010 8602 9010 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 5704 12138 5704 12138 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 5612 18190 5612 18190 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 6670 12750 6670 12750 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 5842 13804 5842 13804 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 8694 12750 8694 12750 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 6256 16014 6256 16014 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 7222 14977 7222 14977 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 8096 13158 8096 13158 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 7314 16150 7314 16150 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 7544 17102 7544 17102 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 8740 18598 8740 18598 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 9062 14382 9062 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 9146 8786 9146 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 14306 7412 14306 7412 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 8234 14416 8234 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9062 15776 9062 15776 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10442 15130 10442 15130 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11868 14042 11868 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8326 11016 8326 11016 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8786 14858 8786 14858 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8970 8058 8970 8058 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8096 8942 8096 8942 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7820 11254 7820 11254 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4140 14042 4140 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4876 11866 4876 11866 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 10810 7344 10810 7344 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4462 14382 4462 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6854 16796 6854 16796 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7038 15402 7038 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8602 12954 8602 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5014 13974 5014 13974 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6026 14042 6026 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 6302 11798 6302 11798 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 5474 12614 5474 12614 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 4922 11730 4922 11730 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 5612 15538 5612 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9982 13158 9982 13158 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 10902 7412 10902 7412 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4784 15402 4784 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7406 15062 7406 15062 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7314 14416 7314 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9384 12206 9384 12206 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 8602 14297 8602 14297 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6946 14008 6946 14008 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10304 13226 10304 13226 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 10810 13481 10810 13481 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8694 14042 8694 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 8096 17714 8096 17714 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10488 17850 10488 17850 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal3 6969 19380 6969 19380 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 7682 17646 7682 17646 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6302 17306 6302 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7544 15674 7544 15674 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10396 14382 10396 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7774 17850 7774 17850 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6808 17034 6808 17034 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10074 14586 10074 14586 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 14398 19040 14398 19040 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6118 19482 6118 19482 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 17020 5610 17020 5610 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 23362 4590 23362 4590 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 20562 4012 20562 4012 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal2 28842 4964 28842 4964 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 22494 6596 22494 6596 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 22557 5202 22557 5202 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 18124 3026 18124 3026 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal2 27186 5474 27186 5474 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23598 6970 23598 6970 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel via1 22143 5202 22143 5202 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 17066 4284 17066 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 25990 4828 25990 4828 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 22527 6290 22527 6290 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 15226 6052 15226 6052 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal2 24886 5916 24886 5916 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 2990 2414 2990 2414 0 ccff_head
rlabel metal2 48622 24694 48622 24694 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2254 24524 2254 24524 0 ccff_tail_0
rlabel metal3 2016 1564 2016 1564 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6222 1472 6222 0 chanx_left_in[11]
rlabel metal3 1004 6460 1004 6460 0 chanx_left_in[12]
rlabel metal1 3082 6902 3082 6902 0 chanx_left_in[13]
rlabel metal1 2990 6290 2990 6290 0 chanx_left_in[14]
rlabel metal2 3726 7531 3726 7531 0 chanx_left_in[15]
rlabel metal2 2438 7429 2438 7429 0 chanx_left_in[16]
rlabel metal1 2990 7854 2990 7854 0 chanx_left_in[17]
rlabel metal2 1794 7837 1794 7837 0 chanx_left_in[18]
rlabel metal1 2484 7378 2484 7378 0 chanx_left_in[19]
rlabel metal3 1740 1972 1740 1972 0 chanx_left_in[1]
rlabel metal2 1610 9673 1610 9673 0 chanx_left_in[20]
rlabel metal1 2990 8942 2990 8942 0 chanx_left_in[21]
rlabel metal1 2599 7854 2599 7854 0 chanx_left_in[22]
rlabel metal2 2806 9707 2806 9707 0 chanx_left_in[23]
rlabel metal3 1717 11356 1717 11356 0 chanx_left_in[24]
rlabel metal2 1610 10931 1610 10931 0 chanx_left_in[25]
rlabel metal1 1472 12206 1472 12206 0 chanx_left_in[26]
rlabel metal3 1188 12580 1188 12580 0 chanx_left_in[27]
rlabel metal1 1794 7820 1794 7820 0 chanx_left_in[28]
rlabel metal1 1472 12818 1472 12818 0 chanx_left_in[29]
rlabel metal1 2576 2482 2576 2482 0 chanx_left_in[2]
rlabel metal1 1472 2958 1472 2958 0 chanx_left_in[3]
rlabel metal1 1472 3502 1472 3502 0 chanx_left_in[4]
rlabel metal3 1004 3604 1004 3604 0 chanx_left_in[5]
rlabel metal1 2990 4114 2990 4114 0 chanx_left_in[6]
rlabel metal2 1794 4267 1794 4267 0 chanx_left_in[7]
rlabel metal1 1472 4658 1472 4658 0 chanx_left_in[8]
rlabel metal1 1472 5202 1472 5202 0 chanx_left_in[9]
rlabel metal2 2806 13583 2806 13583 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal2 2806 18819 2806 18819 0 chanx_left_out[11]
rlabel metal2 2898 19227 2898 19227 0 chanx_left_out[12]
rlabel metal3 1694 19108 1694 19108 0 chanx_left_out[13]
rlabel metal2 2990 19720 2990 19720 0 chanx_left_out[14]
rlabel metal3 1050 19924 1050 19924 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 3266 22015 3266 22015 0 chanx_left_out[20]
rlabel metal3 1487 22372 1487 22372 0 chanx_left_out[21]
rlabel metal1 5474 20502 5474 20502 0 chanx_left_out[22]
rlabel metal1 7222 19414 7222 19414 0 chanx_left_out[23]
rlabel metal1 8096 21862 8096 21862 0 chanx_left_out[24]
rlabel metal2 5060 20196 5060 20196 0 chanx_left_out[25]
rlabel metal2 5244 19924 5244 19924 0 chanx_left_out[26]
rlabel metal1 6532 18190 6532 18190 0 chanx_left_out[27]
rlabel metal2 7544 20740 7544 20740 0 chanx_left_out[28]
rlabel metal1 3864 16150 3864 16150 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel metal1 5290 8534 5290 8534 0 chany_top_in[0]
rlabel metal1 34638 22406 34638 22406 0 chany_top_in[10]
rlabel metal1 32269 24310 32269 24310 0 chany_top_in[11]
rlabel metal2 30130 25041 30130 25041 0 chany_top_in[12]
rlabel metal1 31050 24174 31050 24174 0 chany_top_in[13]
rlabel metal2 35742 22780 35742 22780 0 chany_top_in[14]
rlabel metal1 32200 24174 32200 24174 0 chany_top_in[15]
rlabel metal2 36294 23494 36294 23494 0 chany_top_in[16]
rlabel metal2 33350 24412 33350 24412 0 chany_top_in[17]
rlabel metal2 34086 25245 34086 25245 0 chany_top_in[18]
rlabel metal1 34776 24174 34776 24174 0 chany_top_in[19]
rlabel metal2 27830 23834 27830 23834 0 chany_top_in[1]
rlabel metal1 36018 24072 36018 24072 0 chany_top_in[20]
rlabel metal1 36708 24174 36708 24174 0 chany_top_in[21]
rlabel metal1 36662 23698 36662 23698 0 chany_top_in[22]
rlabel metal1 37490 24174 37490 24174 0 chany_top_in[23]
rlabel metal1 37812 23698 37812 23698 0 chany_top_in[24]
rlabel metal2 38502 25245 38502 25245 0 chany_top_in[25]
rlabel metal2 39238 25245 39238 25245 0 chany_top_in[26]
rlabel metal1 39836 24242 39836 24242 0 chany_top_in[27]
rlabel metal1 41078 24174 41078 24174 0 chany_top_in[28]
rlabel metal1 41354 23698 41354 23698 0 chany_top_in[29]
rlabel metal3 17204 22168 17204 22168 0 chany_top_in[2]
rlabel metal3 17204 22440 17204 22440 0 chany_top_in[3]
rlabel metal2 14490 23681 14490 23681 0 chany_top_in[4]
rlabel metal1 17204 22746 17204 22746 0 chany_top_in[5]
rlabel metal2 29210 24225 29210 24225 0 chany_top_in[6]
rlabel metal1 28566 24140 28566 24140 0 chany_top_in[7]
rlabel metal1 29578 23664 29578 23664 0 chany_top_in[8]
rlabel metal1 31372 23698 31372 23698 0 chany_top_in[9]
rlabel metal1 3634 23154 3634 23154 0 chany_top_out[0]
rlabel metal1 8234 24276 8234 24276 0 chany_top_out[10]
rlabel metal1 9568 23766 9568 23766 0 chany_top_out[11]
rlabel metal2 10718 24497 10718 24497 0 chany_top_out[12]
rlabel metal2 11270 24184 11270 24184 0 chany_top_out[13]
rlabel metal2 12558 21556 12558 21556 0 chany_top_out[14]
rlabel metal2 12558 25034 12558 25034 0 chany_top_out[15]
rlabel metal2 13301 26316 13301 26316 0 chany_top_out[16]
rlabel metal2 13846 25204 13846 25204 0 chany_top_out[17]
rlabel metal1 13570 24276 13570 24276 0 chany_top_out[18]
rlabel metal1 15364 22202 15364 22202 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 14996 23766 14996 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal2 17211 26316 17211 26316 0 chany_top_out[22]
rlabel metal1 16974 23154 16974 23154 0 chany_top_out[23]
rlabel metal1 17250 23766 17250 23766 0 chany_top_out[24]
rlabel metal1 16468 24242 16468 24242 0 chany_top_out[25]
rlabel metal2 17894 23460 17894 23460 0 chany_top_out[26]
rlabel metal1 20930 22100 20930 22100 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal2 21574 25272 21574 25272 0 chany_top_out[29]
rlabel metal1 4094 23766 4094 23766 0 chany_top_out[2]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7360 21930 7360 21930 0 chany_top_out[6]
rlabel metal1 6486 24242 6486 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8694 24422 8694 24422 0 chany_top_out[9]
rlabel metal2 18446 17408 18446 17408 0 clknet_0_prog_clk
rlabel metal1 7498 10506 7498 10506 0 clknet_4_0_0_prog_clk
rlabel metal1 22310 11662 22310 11662 0 clknet_4_10_0_prog_clk
rlabel metal2 22034 16320 22034 16320 0 clknet_4_11_0_prog_clk
rlabel metal1 19734 19244 19734 19244 0 clknet_4_12_0_prog_clk
rlabel metal1 19734 20502 19734 20502 0 clknet_4_13_0_prog_clk
rlabel metal1 27968 18258 27968 18258 0 clknet_4_14_0_prog_clk
rlabel metal2 37858 22882 37858 22882 0 clknet_4_15_0_prog_clk
rlabel metal1 8372 12614 8372 12614 0 clknet_4_1_0_prog_clk
rlabel metal1 14536 10030 14536 10030 0 clknet_4_2_0_prog_clk
rlabel metal2 14306 13090 14306 13090 0 clknet_4_3_0_prog_clk
rlabel metal1 4554 17646 4554 17646 0 clknet_4_4_0_prog_clk
rlabel metal2 9430 19040 9430 19040 0 clknet_4_5_0_prog_clk
rlabel metal2 14582 19652 14582 19652 0 clknet_4_6_0_prog_clk
rlabel metal1 12788 21522 12788 21522 0 clknet_4_7_0_prog_clk
rlabel metal2 16882 7616 16882 7616 0 clknet_4_8_0_prog_clk
rlabel metal1 19964 12750 19964 12750 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25576 2414 25576 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28382 1581 28382 1581 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33580 2414 33580 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 14766 1622 14766 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17434 1622 17434 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 20102 959 20102 959 0 gfpga_pad_io_soc_out[2]
rlabel metal2 22770 1622 22770 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal1 5060 2618 5060 2618 0 net1
rlabel metal2 8970 15997 8970 15997 0 net10
rlabel metal1 10787 16966 10787 16966 0 net100
rlabel metal1 4002 16490 4002 16490 0 net101
rlabel metal2 19458 19839 19458 19839 0 net102
rlabel metal1 8648 19346 8648 19346 0 net103
rlabel metal2 3542 15606 3542 15606 0 net104
rlabel metal1 2277 14382 2277 14382 0 net105
rlabel metal1 1794 15028 1794 15028 0 net106
rlabel metal2 3450 14756 3450 14756 0 net107
rlabel metal1 2277 16082 2277 16082 0 net108
rlabel metal1 2760 16558 2760 16558 0 net109
rlabel metal1 11546 16626 11546 16626 0 net11
rlabel metal2 1794 17255 1794 17255 0 net110
rlabel metal1 1794 17680 1794 17680 0 net111
rlabel metal1 1794 18292 1794 18292 0 net112
rlabel metal2 2254 15538 2254 15538 0 net113
rlabel metal3 4623 9588 4623 9588 0 net114
rlabel metal3 6900 13532 6900 13532 0 net115
rlabel metal2 33626 24718 33626 24718 0 net116
rlabel metal2 35650 24616 35650 24616 0 net117
rlabel metal2 33810 24174 33810 24174 0 net118
rlabel metal2 31786 23936 31786 23936 0 net119
rlabel metal1 1518 6630 1518 6630 0 net12
rlabel metal2 32062 24072 32062 24072 0 net120
rlabel metal1 10028 24174 10028 24174 0 net121
rlabel metal2 34822 24514 34822 24514 0 net122
rlabel metal2 33718 24004 33718 24004 0 net123
rlabel metal1 2300 24174 2300 24174 0 net124
rlabel metal2 13202 20604 13202 20604 0 net125
rlabel metal1 15962 22610 15962 22610 0 net126
rlabel via3 17043 20740 17043 20740 0 net127
rlabel metal2 15502 22865 15502 22865 0 net128
rlabel metal2 14352 17612 14352 17612 0 net129
rlabel metal1 2162 7514 2162 7514 0 net13
rlabel metal2 17342 20468 17342 20468 0 net130
rlabel metal2 33902 23171 33902 23171 0 net131
rlabel metal2 20378 22039 20378 22039 0 net132
rlabel metal1 19320 20026 19320 20026 0 net133
rlabel metal2 22034 24480 22034 24480 0 net134
rlabel metal2 3864 17204 3864 17204 0 net135
rlabel metal1 14122 22440 14122 22440 0 net136
rlabel metal2 15134 23613 15134 23613 0 net137
rlabel metal2 2438 16558 2438 16558 0 net138
rlabel metal1 7084 21998 7084 21998 0 net139
rlabel metal2 12650 5916 12650 5916 0 net14
rlabel metal2 2024 18292 2024 18292 0 net140
rlabel metal3 6233 20740 6233 20740 0 net141
rlabel metal3 5221 19380 5221 19380 0 net142
rlabel metal1 4968 2414 4968 2414 0 net143
rlabel metal1 7682 2414 7682 2414 0 net144
rlabel metal1 9706 2414 9706 2414 0 net145
rlabel metal1 12420 2414 12420 2414 0 net146
rlabel metal2 15042 3162 15042 3162 0 net147
rlabel metal1 17204 2822 17204 2822 0 net148
rlabel metal1 19136 2822 19136 2822 0 net149
rlabel metal2 12098 18564 12098 18564 0 net15
rlabel metal1 22356 2414 22356 2414 0 net150
rlabel metal1 21850 21522 21850 21522 0 net151
rlabel metal2 23414 20706 23414 20706 0 net152
rlabel metal2 17618 18972 17618 18972 0 net153
rlabel metal1 23828 21930 23828 21930 0 net154
rlabel metal1 23092 22746 23092 22746 0 net155
rlabel metal1 24610 23834 24610 23834 0 net156
rlabel metal1 27646 22066 27646 22066 0 net157
rlabel metal1 26358 19482 26358 19482 0 net158
rlabel metal1 28658 18394 28658 18394 0 net159
rlabel metal2 5750 15929 5750 15929 0 net16
rlabel metal2 14674 19380 14674 19380 0 net160
rlabel metal1 20378 17578 20378 17578 0 net161
rlabel metal1 24150 18802 24150 18802 0 net162
rlabel metal1 12512 20366 12512 20366 0 net163
rlabel metal2 20470 16830 20470 16830 0 net164
rlabel metal1 14122 8874 14122 8874 0 net165
rlabel metal1 14168 8466 14168 8466 0 net166
rlabel metal1 10580 6834 10580 6834 0 net167
rlabel metal2 11914 8194 11914 8194 0 net168
rlabel metal2 13570 12002 13570 12002 0 net169
rlabel metal1 4186 7718 4186 7718 0 net17
rlabel metal1 13432 7514 13432 7514 0 net170
rlabel metal1 17020 16626 17020 16626 0 net171
rlabel metal2 15410 17034 15410 17034 0 net172
rlabel metal1 14996 15470 14996 15470 0 net173
rlabel metal1 8418 11866 8418 11866 0 net174
rlabel metal2 9430 10030 9430 10030 0 net175
rlabel metal2 8694 15521 8694 15521 0 net176
rlabel metal1 12144 18258 12144 18258 0 net177
rlabel metal1 20700 14926 20700 14926 0 net178
rlabel metal2 9246 20043 9246 20043 0 net179
rlabel metal1 8234 16558 8234 16558 0 net18
rlabel metal2 4692 17204 4692 17204 0 net180
rlabel metal2 12558 8704 12558 8704 0 net181
rlabel metal1 5934 9622 5934 9622 0 net182
rlabel metal1 32936 23834 32936 23834 0 net183
rlabel via2 9798 21301 9798 21301 0 net184
rlabel metal1 10672 18258 10672 18258 0 net185
rlabel metal2 14122 14756 14122 14756 0 net186
rlabel metal1 10626 15402 10626 15402 0 net187
rlabel metal1 16054 12750 16054 12750 0 net188
rlabel metal1 16146 8602 16146 8602 0 net189
rlabel metal1 13478 16694 13478 16694 0 net19
rlabel metal1 7452 10778 7452 10778 0 net190
rlabel metal1 5750 12886 5750 12886 0 net191
rlabel metal1 15594 13158 15594 13158 0 net192
rlabel metal2 12466 14161 12466 14161 0 net193
rlabel metal1 27968 16558 27968 16558 0 net194
rlabel via2 32154 23579 32154 23579 0 net195
rlabel metal2 36018 23953 36018 23953 0 net196
rlabel metal1 18676 16558 18676 16558 0 net197
rlabel metal1 16422 20774 16422 20774 0 net198
rlabel metal2 48438 22746 48438 22746 0 net2
rlabel metal2 3404 15980 3404 15980 0 net20
rlabel metal1 6946 16626 6946 16626 0 net21
rlabel metal1 2070 11662 2070 11662 0 net22
rlabel metal2 2530 13129 2530 13129 0 net23
rlabel metal2 1886 12954 1886 12954 0 net24
rlabel metal1 3404 2346 3404 2346 0 net25
rlabel metal1 1886 3060 1886 3060 0 net26
rlabel via1 13202 8891 13202 8891 0 net27
rlabel metal2 13386 8092 13386 8092 0 net28
rlabel metal2 10626 6256 10626 6256 0 net29
rlabel metal1 7176 3706 7176 3706 0 net3
rlabel metal2 9706 6358 9706 6358 0 net30
rlabel metal2 11822 14654 11822 14654 0 net31
rlabel metal1 5888 5134 5888 5134 0 net32
rlabel metal1 16882 19686 16882 19686 0 net33
rlabel metal2 34546 23001 34546 23001 0 net34
rlabel metal1 11684 16422 11684 16422 0 net35
rlabel metal2 12466 16813 12466 16813 0 net36
rlabel metal1 28106 20570 28106 20570 0 net37
rlabel metal2 35558 22304 35558 22304 0 net38
rlabel metal2 31878 23834 31878 23834 0 net39
rlabel metal1 14168 14042 14168 14042 0 net4
rlabel metal2 36110 23086 36110 23086 0 net40
rlabel metal2 33534 24565 33534 24565 0 net41
rlabel metal2 34270 24820 34270 24820 0 net42
rlabel metal2 34638 24548 34638 24548 0 net43
rlabel via2 17434 20893 17434 20893 0 net44
rlabel metal1 13294 15674 13294 15674 0 net45
rlabel metal1 36294 24038 36294 24038 0 net46
rlabel metal2 36754 22542 36754 22542 0 net47
rlabel metal2 37490 23936 37490 23936 0 net48
rlabel metal1 36248 23562 36248 23562 0 net49
rlabel metal2 13294 12716 13294 12716 0 net5
rlabel via2 16974 15861 16974 15861 0 net50
rlabel metal1 16422 19482 16422 19482 0 net51
rlabel metal2 40342 24412 40342 24412 0 net52
rlabel metal2 41354 24089 41354 24089 0 net53
rlabel metal1 41354 23596 41354 23596 0 net54
rlabel metal1 23644 20774 23644 20774 0 net55
rlabel metal1 19044 20570 19044 20570 0 net56
rlabel metal2 14306 24548 14306 24548 0 net57
rlabel metal1 26496 24174 26496 24174 0 net58
rlabel metal1 25484 22950 25484 22950 0 net59
rlabel metal1 2898 6664 2898 6664 0 net6
rlabel metal1 26772 23018 26772 23018 0 net60
rlabel metal1 27140 22746 27140 22746 0 net61
rlabel metal1 14720 21998 14720 21998 0 net62
rlabel metal2 25530 4114 25530 4114 0 net63
rlabel metal1 25806 4522 25806 4522 0 net64
rlabel metal1 29808 2618 29808 2618 0 net65
rlabel metal2 33534 3842 33534 3842 0 net66
rlabel metal1 27462 5610 27462 5610 0 net67
rlabel metal1 40020 22746 40020 22746 0 net68
rlabel metal2 44022 21437 44022 21437 0 net69
rlabel metal1 5980 7174 5980 7174 0 net7
rlabel metal2 41630 20944 41630 20944 0 net70
rlabel metal2 46874 22253 46874 22253 0 net71
rlabel metal2 46966 22576 46966 22576 0 net72
rlabel metal2 45310 20604 45310 20604 0 net73
rlabel metal2 48714 19720 48714 19720 0 net74
rlabel metal2 41446 20774 41446 20774 0 net75
rlabel metal2 44482 21369 44482 21369 0 net76
rlabel metal2 48346 20944 48346 20944 0 net77
rlabel metal2 48806 19958 48806 19958 0 net78
rlabel metal2 49266 19414 49266 19414 0 net79
rlabel metal1 7958 15402 7958 15402 0 net8
rlabel metal2 48530 22440 48530 22440 0 net80
rlabel metal1 47794 21318 47794 21318 0 net81
rlabel metal1 6578 19278 6578 19278 0 net82
rlabel metal1 1794 13260 1794 13260 0 net83
rlabel metal1 13386 19176 13386 19176 0 net84
rlabel metal1 1794 19380 1794 19380 0 net85
rlabel metal1 1794 19924 1794 19924 0 net86
rlabel metal2 1794 21964 1794 21964 0 net87
rlabel metal1 1840 20910 1840 20910 0 net88
rlabel metal1 1794 21590 1794 21590 0 net89
rlabel metal1 7728 14926 7728 14926 0 net9
rlabel metal1 3864 20434 3864 20434 0 net90
rlabel metal1 2898 21998 2898 21998 0 net91
rlabel metal1 1840 22610 1840 22610 0 net92
rlabel metal1 1886 23086 1886 23086 0 net93
rlabel via2 1794 13923 1794 13923 0 net94
rlabel metal1 4416 21998 4416 21998 0 net95
rlabel metal1 3680 19346 3680 19346 0 net96
rlabel metal2 6118 21148 6118 21148 0 net97
rlabel metal3 4186 16660 4186 16660 0 net98
rlabel metal1 6118 12682 6118 12682 0 net99
rlabel metal2 38778 2098 38778 2098 0 prog_clk
rlabel metal1 41860 24378 41860 24378 0 prog_reset_top_in
rlabel metal1 18446 16966 18446 16966 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal1 25760 19890 25760 19890 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal1 29900 16626 29900 16626 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 13524 20366 13524 20366 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal1 17204 23018 17204 23018 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal1 18722 22474 18722 22474 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 18492 22542 18492 22542 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal1 19044 23766 19044 23766 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal2 15134 21250 15134 21250 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal1 21850 22746 21850 22746 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal2 20470 20825 20470 20825 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal1 24104 23562 24104 23562 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 23920 21454 23920 21454 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 23828 21590 23828 21590 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal1 26450 18938 26450 18938 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 26910 20366 26910 20366 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 18584 19890 18584 19890 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 20509 19142 20509 19142 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 26266 22066 26266 22066 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal2 27646 20366 27646 20366 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal1 26450 23494 26450 23494 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal1 27738 22576 27738 22576 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal2 29026 23936 29026 23936 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal1 28842 23494 28842 23494 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal1 28658 21454 28658 21454 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal1 31142 22134 31142 22134 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 27462 19414 27462 19414 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal1 29578 21318 29578 21318 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 28612 18054 28612 18054 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 29348 19142 29348 19142 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 20102 19890 20102 19890 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal2 19734 21148 19734 21148 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 28842 17408 28842 17408 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 20654 19822 20654 19822 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 21758 19686 21758 19686 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 19090 20400 19090 20400 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 25070 15062 25070 15062 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal1 37743 22406 37743 22406 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal2 25162 16065 25162 16065 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 20654 13804 20654 13804 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 17250 9962 17250 9962 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal2 24058 11968 24058 11968 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 21436 12750 21436 12750 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 16284 8874 16284 8874 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 20194 14450 20194 14450 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 15548 10098 15548 10098 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal1 14674 9486 14674 9486 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 16008 12274 16008 12274 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal2 15042 9928 15042 9928 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 17434 13668 17434 13668 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 16882 13226 16882 13226 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 21206 9690 21206 9690 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 22724 11798 22724 11798 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 24150 10744 24150 10744 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 18124 15334 18124 15334 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal2 17342 14722 17342 14722 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal2 16330 14620 16330 14620 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 14996 15062 14996 15062 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15548 13498 15548 13498 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal1 15502 13362 15502 13362 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal2 11546 10370 11546 10370 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal2 12098 11798 12098 11798 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 12972 9350 12972 9350 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal2 12006 9860 12006 9860 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12282 13906 12282 13906 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 12328 12274 12328 12274 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12282 17136 12282 17136 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal2 13754 14722 13754 14722 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 13478 19788 13478 19788 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal1 13570 17850 13570 17850 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal2 9062 20060 9062 20060 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal1 11730 20366 11730 20366 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 4876 18666 4876 18666 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 8096 16014 8096 16014 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 19826 13226 19826 13226 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal1 22770 11322 22770 11322 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 17066 9486 17066 9486 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 7912 21590 7912 21590 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal1 7406 18598 7406 18598 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 10304 22950 10304 22950 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal1 9430 21624 9430 21624 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13386 21624 13386 21624 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal1 13386 22950 13386 22950 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 15180 19890 15180 19890 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal2 14030 20196 14030 20196 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 16790 17714 16790 17714 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal2 20102 18428 20102 18428 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 18492 17102 18492 17102 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 21942 14824 21942 14824 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal1 21390 17068 21390 17068 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 20240 15402 20240 15402 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 24196 14246 24196 14246 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 20378 10336 20378 10336 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal2 14858 18632 14858 18632 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 25162 19958 25162 19958 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27278 16422 27278 16422 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21114 19006 21114 19006 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4324 12886 4324 12886 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 12374 24242 12374 24242 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 8119 12444 8119 12444 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 26634 18275 26634 18275 0 sb_8__0_.mux_left_track_13.out
rlabel metal1 16882 21658 16882 21658 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 15594 21403 15594 21403 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6440 21998 6440 21998 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 15594 20910 15594 20910 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16514 20655 16514 20655 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3680 12818 3680 12818 0 sb_8__0_.mux_left_track_17.out
rlabel metal1 24794 23086 24794 23086 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 15847 20740 15847 20740 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 15368 19458 15368 0 sb_8__0_.mux_left_track_19.out
rlabel metal1 23000 21658 23000 21658 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 15674 19642 15674 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7728 15062 7728 15062 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 24886 20230 24886 20230 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 10718 12835 10718 12835 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31970 18105 31970 18105 0 sb_8__0_.mux_left_track_3.out
rlabel metal1 18032 19822 18032 19822 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 20179 17250 20179 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16146 17510 16146 17510 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 27324 21658 27324 21658 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20378 21369 20378 21369 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2392 23698 2392 23698 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 24610 21998 24610 21998 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22310 11327 22310 11327 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 9200 13668 9200 13668 0 sb_8__0_.mux_left_track_35.out
rlabel metal1 30498 22406 30498 22406 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23736 17238 23736 17238 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 15997 21298 15997 0 sb_8__0_.mux_left_track_45.out
rlabel metal1 30130 21896 30130 21896 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24978 21318 24978 21318 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12190 16048 12190 16048 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 25208 20978 25208 20978 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23966 18224 23966 18224 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 13110 15147 13110 15147 0 sb_8__0_.mux_left_track_49.out
rlabel metal2 30222 19516 30222 19516 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21574 16456 21574 16456 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17250 21862 17250 21862 0 sb_8__0_.mux_left_track_5.out
rlabel metal1 17250 20570 17250 20570 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16928 20230 16928 20230 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5750 13719 5750 13719 0 sb_8__0_.mux_left_track_51.out
rlabel metal2 21206 17204 21206 17204 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16974 16082 16974 16082 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13938 18632 13938 18632 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 22586 19414 22586 19414 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 19482 22862 19482 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 18666 14858 18666 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel via3 7107 12852 7107 12852 0 sb_8__0_.mux_left_track_9.out
rlabel metal1 18538 20536 18538 20536 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 19686 13202 19686 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21206 21053 21206 21053 0 sb_8__0_.mux_top_track_0.out
rlabel metal2 27094 17408 27094 17408 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27738 16490 27738 16490 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26634 16456 26634 16456 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23414 19346 23414 19346 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23598 19108 23598 19108 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18906 16082 18906 16082 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 21390 12818 21390 12818 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21160 12954 21160 12954 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 12614 20838 12614 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14536 9078 14536 9078 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal3 17204 14756 17204 14756 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 14398 16473 14398 16473 0 sb_8__0_.mux_top_track_12.out
rlabel metal1 16054 10540 16054 10540 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14858 8602 14858 8602 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14720 16558 14720 16558 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14858 9044 14858 9044 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 15088 10778 15088 10778 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 10608 14766 10608 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14398 10744 14398 10744 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 10994 15963 10994 15963 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 17986 11866 17986 11866 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12673 12818 12673 12818 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11178 14518 11178 14518 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20930 21862 20930 21862 0 sb_8__0_.mux_top_track_18.out
rlabel metal2 17894 16694 17894 16694 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13202 14144 13202 14144 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17388 15946 17388 15946 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19090 19652 19090 19652 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 24840 13974 24840 13974 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25392 14042 25392 14042 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 9622 22080 9622 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 8058 15134 8058 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19182 19346 19182 19346 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33396 22406 33396 22406 0 sb_8__0_.mux_top_track_20.out
rlabel metal2 15870 16354 15870 16354 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11730 15470 11730 15470 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34822 23698 34822 23698 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 14398 13804 14398 13804 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19044 14382 19044 14382 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 9430 13379 9430 13379 0 sb_8__0_.mux_top_track_24.out
rlabel metal1 14168 12614 14168 12614 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13662 14382 13662 14382 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32292 23018 32292 23018 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 10626 11934 10626 11934 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4002 21063 4002 21063 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32660 22610 32660 22610 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 10442 10234 10442 10234 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10856 8942 10856 8942 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 29762 21454 29762 21454 0 sb_8__0_.mux_top_track_30.out
rlabel metal2 12558 13872 12558 13872 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 12098 15589 12098 15589 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33074 23698 33074 23698 0 sb_8__0_.mux_top_track_32.out
rlabel metal1 12834 15130 12834 15130 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 31786 20111 31786 20111 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32384 23630 32384 23630 0 sb_8__0_.mux_top_track_34.out
rlabel metal2 12558 17867 12558 17867 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10442 19431 10442 19431 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1610 11016 1610 11016 0 sb_8__0_.mux_top_track_36.out
rlabel metal2 11546 21964 11546 21964 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 2346 11186 2346 11186 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4738 9554 4738 9554 0 sb_8__0_.mux_top_track_38.out
rlabel metal1 6118 16218 6118 16218 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 5152 20060 5152 20060 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 16422 18814 16422 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 20654 12648 20654 12648 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19182 12954 19182 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17388 12954 17388 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13248 13838 13248 13838 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16422 14042 16422 14042 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5566 8602 5566 8602 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7728 17306 7728 17306 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 6555 10404 6555 10404 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 8194 9154 8194 0 sb_8__0_.mux_top_track_42.out
rlabel metal2 10626 20910 10626 20910 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 8349 20876 8349 20876 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32522 17340 32522 17340 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 16192 19414 16192 19414 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12190 20740 12190 20740 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32430 20655 32430 20655 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32844 21998 32844 21998 0 sb_8__0_.mux_top_track_46.out
rlabel metal1 18262 18870 18262 18870 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12834 18904 12834 18904 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13202 20026 13202 20026 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 2162 10710 2162 10710 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 17526 18122 17526 18122 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14398 17034 14398 17034 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15134 18343 15134 18343 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19458 14739 19458 14739 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 19044 18394 19044 18394 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13662 16422 13662 16422 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 13872 19642 13872 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 32982 22627 32982 22627 0 sb_8__0_.mux_top_track_6.out
rlabel metal2 20746 16830 20746 16830 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 16558 22862 16558 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 15062 20930 15062 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20056 14994 20056 14994 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel via1 19734 14875 19734 14875 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18354 17714 18354 17714 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 23322 13396 23322 13396 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 13226 23276 13226 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21666 13668 21666 13668 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15594 8568 15594 8568 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19872 14042 19872 14042 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 44758 25340 44758 25340 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45494 25296 45494 25296 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46368 24174 46368 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 46736 23698 46736 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48254 24174 48254 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 43378 23834 43378 23834 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 44252 23698 44252 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 49542 22185 49542 22185 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 49358 22831 49358 22831 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 49542 23953 49542 23953 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 48346 24259 48346 24259 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 41446 2948 41446 2948 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 44114 2200 44114 2200 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 27554 4114 27554 4114 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 26542 5576 26542 5576 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
