* NGSPICE file created from top_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

.subckt top_tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ bottom_width_0_height_0_subtile_0__pin_reg_out_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ bottom_width_0_height_0_subtile_2__pin_inpad_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0] chanx_right_in_0[10]
+ chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13] chanx_right_in_0[14]
+ chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17] chanx_right_in_0[18]
+ chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20] chanx_right_in_0[21]
+ chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24] chanx_right_in_0[25]
+ chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28] chanx_right_in_0[29]
+ chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4] chanx_right_in_0[5]
+ chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8] chanx_right_in_0[9]
+ chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11] chanx_right_out_0[12]
+ chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15] chanx_right_out_0[16]
+ chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19] chanx_right_out_0[1]
+ chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22] chanx_right_out_0[23]
+ chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26] chanx_right_out_0[27]
+ chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2] chanx_right_out_0[3]
+ chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6] chanx_right_out_0[7]
+ chanx_right_out_0[8] chanx_right_out_0[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] clk0 gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk
+ prog_reset reset right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
+ right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ right_width_0_height_0_subtile_0__pin_O_10_ right_width_0_height_0_subtile_0__pin_O_11_
+ right_width_0_height_0_subtile_0__pin_O_12_ right_width_0_height_0_subtile_0__pin_O_13_
+ right_width_0_height_0_subtile_0__pin_O_14_ right_width_0_height_0_subtile_0__pin_O_15_
+ right_width_0_height_0_subtile_0__pin_O_8_ right_width_0_height_0_subtile_0__pin_O_9_
+ sc_in sc_out test_enable top_width_0_height_0_subtile_0__pin_O_0_ top_width_0_height_0_subtile_0__pin_O_1_
+ top_width_0_height_0_subtile_0__pin_O_2_ top_width_0_height_0_subtile_0__pin_O_3_
+ top_width_0_height_0_subtile_0__pin_O_4_ top_width_0_height_0_subtile_0__pin_O_5_
+ top_width_0_height_0_subtile_0__pin_O_6_ top_width_0_height_0_subtile_0__pin_O_7_
+ top_width_0_height_0_subtile_0__pin_cin_0_ top_width_0_height_0_subtile_0__pin_reg_in_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.out sky130_fd_sc_hd__buf_4
XFILLER_89_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_3__S sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_11.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_294_ net14 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input92_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_1__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__304__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_1_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_346_ sb_1__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_277_ net38 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_3__261 VGND VGND VPWR VPWR net261 cby_1__8_.mux_right_ipin_4.mux_l2_in_3__261/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput231 net231 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
Xoutput220 net220 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_15_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_2.mem_out\[2\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_12.mux_l3_in_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input55_A chanx_right_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_1_ net6 cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_329_ sb_1__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_13.mux_l3_in_0_ sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_4.mux_l2_in_3__359 VGND VGND VPWR VPWR net359 sb_1__8_.mux_right_track_4.mux_l2_in_3__359/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk
+ sb_1__8_.mem_bottom_track_33.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_35.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1__A0 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__312__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l1_in_2__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__365 VGND VGND VPWR VPWR net365
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__365/LO sky130_fd_sc_hd__conb_1
XFILLER_13_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_1_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_52.mux_l1_in_1__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__241 VGND VGND VPWR VPWR net241 cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__241/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2_ net43 net12 cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_12.mux_l1_in_3_ net354 net26 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_39_prog_clk sb_1__8_.mem_right_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_3__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_13.mux_l2_in_1_ net317 net6 sb_1__8_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__307__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_11.mux_l2_in_3__342 VGND VGND VPWR VPWR net342 sb_1__8_.mux_left_track_11.mux_l2_in_3__342/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_1.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_44.mux_l1_in_1__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_3.mux_l1_in_1__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_6.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_1__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk sb_1__8_.mem_left_track_11.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_85_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_10.mux_l2_in_3__353 VGND VGND VPWR VPWR net353 sb_1__8_.mux_right_track_10.mux_l2_in_3__353/LO
+ sky130_fd_sc_hd__conb_1
X_362_ net117 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ sb_1__8_.mux_left_track_1.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input85_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2__A0 net29 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__314
+ VGND VGND VPWR VPWR net314 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__314/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__369 VGND VGND VPWR VPWR net369 cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__369/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_11.mux_l2_in_3__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_12.mux_l3_in_0_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_3.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2__A1 net41 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out
+ net18 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__268
+ VGND VGND VPWR VPWR net268 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__268/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_345_ sb_1__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net308 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_2__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_276_ net37 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__315__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput210 net210 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput232 net232 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_15_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_2.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__A1 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A chanx_right_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_12.mux_l2_in_1_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_328_ sb_1__8_.mux_bottom_track_51.out VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_load_slew238_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net297 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_11.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input102_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_bottom_track_11.mux_l1_in_1__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_52.mux_l1_in_1__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net268 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_12.mux_l1_in_2_ net12 net86 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk sb_1__8_.mem_right_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_0__S sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_13.mux_l2_in_0_ net11 sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_2__S sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net270 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__mux2_4
Xcby_1__8_.mux_right_ipin_1.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_15_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND
+ VPWR VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_3.mux_l1_in_1__A1 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_1__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_3__256 VGND VGND VPWR VPWR net256 cby_1__8_.mux_right_ipin_13.mux_l2_in_3__256/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk sb_1__8_.mem_left_track_11.ccff_head
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_85_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_2__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_361_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ sb_1__8_.mux_left_track_3.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input78_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2__A1 net37 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output234_A net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_3.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_43.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out
+ net21 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_14.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_2__A0 sb_1__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_0.mux_l2_in_3_ net352 net4 sb_1__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
X_344_ sb_1__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_2__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_275_ sb_1__8_.mux_left_track_37.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput200 net200 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
XANTENNA_cby_1__8_.mux_right_ipin_1.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput211 net211 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
XANTENNA__331__A sb_1__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_2.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_28_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__291
+ VGND VGND VPWR VPWR net291 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__291/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1__A0 sb_1__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_12.mux_l2_in_0_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_327_ net52 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_3__S sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__326__A net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_bottom_track_11.mux_l1_in_1__A1 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input60_A chanx_right_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk sb_1__8_.mem_right_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l2_in_2__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_7.mux_l2_in_3_ net351 net233 sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_0.mux_l4_in_0_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sb_1__8_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_25_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_12.mux_l1_in_1_ net68 net80 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_11.mux_l2_in_3__A1 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_right_track_0.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_3.mux_l1_in_0__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND
+ VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput100 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_49.mux_l1_in_0__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_0.mux_l3_in_1_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net114 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net299 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__mux2_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_2__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_360_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_291_ sb_1__8_.mux_left_track_5.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net119 net97 VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_13.mux_l1_in_0_ net224 net41 sb_1__8_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_7.mux_l4_in_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output227_A net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ sb_1__8_.mem_bottom_track_21.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_21.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_25.mux_l2_in_0_ sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_25.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__329__A sb_1__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_3.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_23_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_37.mux_l3_in_0_ sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out
+ net24 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_0.mux_l2_in_2_ net21 net92 sb_1__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ sb_1__8_.mux_bottom_track_21.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input90_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ net35 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput201 net201 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
Xoutput234 net234 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk
+ cbx_1__8_.cbx_1__8_.ccff_head net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_1__8_.mem_right_track_0.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_41.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_7.mux_l3_in_1_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_1__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_25.mux_l1_in_1_ net323 net32 sb_1__8_.mem_bottom_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_7.mux_l1_in_0__A0 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_326_ net53 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__243 VGND VGND VPWR VPWR net243 cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__243/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_37.mux_l2_in_1_ net330 net14 sb_1__8_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_2.mux_l2_in_3__355 VGND VGND VPWR VPWR net355 sb_1__8_.mux_right_track_2.mux_l2_in_3__355/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_13.mux_l1_in_3__343 VGND VGND VPWR VPWR net343 sb_1__8_.mux_left_track_13.mux_l1_in_3__343/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input53_A chanx_right_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_3.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_309_ sb_1__8_.mux_right_track_28.out VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net289 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_7.mux_l2_in_2_ net231 net229 sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_2__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_12.mux_l1_in_0_ net102 net108 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net286 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l2_in_3__A1 sb_1__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_12.mux_l1_in_3__354 VGND VGND VPWR VPWR net354 sb_1__8_.mux_right_track_12.mux_l1_in_3__354/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk cbx_1__8_.cbx_1__8_.ccff_tail net236 VGND VGND VPWR VPWR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_36.mux_l3_in_0_ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_1__A0 sb_1__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_3.mux_l1_in_0__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__277
+ VGND VGND VPWR VPWR net277 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__277/LO
+ sky130_fd_sc_hd__conb_1
Xinput101 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__A0 sb_1__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput112 sc_in VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_7.mux_l1_in_3_ net227 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_1__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_0.mux_l3_in_0_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_1__S sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_39.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__350__A sb_1__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_15.mux_l1_in_0__A0 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_1.mux_l3_in_0_ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_290_ sb_1__8_.mux_left_track_7.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__A0 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2__A0 sb_1__8_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk
+ sb_1__8_.mem_bottom_track_19.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_36.mux_l2_in_1_ net358 sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_1.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__345__A sb_1__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.out sky130_fd_sc_hd__clkbuf_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_0.mux_l2_in_1_ net75 net105 sb_1__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_342_ sb_1__8_.mux_bottom_track_23.out VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_273_ net34 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input83_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l2_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_1.mux_l2_in_1_ net315 sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4__A0 sb_1__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput213 net213 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
Xoutput202 net202 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail net97 VGND
+ VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_7.mux_l3_in_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_1__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_36.mux_l1_in_2_ net8 net89 sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_25.mux_l1_in_0_ net222 net62 sb_1__8_.mem_bottom_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_46_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_7.mux_l1_in_0__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_325_ net54 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_29.mux_l1_in_3_ net345 net231 sb_1__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_37.mux_l2_in_0_ net224 sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_27.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_27.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk cby_1__8_.mem_right_ipin_10.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_95_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input46_A chanx_right_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_1.mux_l1_in_2_ net21 net23 sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ net9 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3_ net371 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_load_slew236_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_7.mux_l2_in_1_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_2__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__8_.mem_right_track_44.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__353__A sb_1__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_2__S sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input100_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__A1 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_23.mux_l1_in_0__A0 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_29.mux_l3_in_0_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xinput102 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net102 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_5.mux_l2_in_1__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput113 test_enable VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_8
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4_ sb_1__8_.mux_left_track_45.out net30
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_3_ net259 net52 cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_7.mux_l1_in_2_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net88 sb_1__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l1_in_2__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__294
+ VGND VGND VPWR VPWR net294 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__294/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_50_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk sb_1__8_.mem_bottom_track_9.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__A0 sb_1__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_15.mux_l1_in_0__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_21.mux_l1_in_1__321 VGND VGND VPWR VPWR net321 sb_1__8_.mux_bottom_track_21.mux_l1_in_1__321/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_3__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3_ net244 sb_1__8_.mux_left_track_45.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_right_track_36.mux_l2_in_0_ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net281 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__mux2_4
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.out sky130_fd_sc_hd__clkbuf_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_10.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_29.mux_l2_in_1_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_90_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_4_ sb_1__8_.mux_bottom_track_41.out net92 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4__A0 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk cby_1__8_.mem_right_ipin_13.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_right_track_0.mux_l2_in_0_ net102 sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_right_track_0.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_341_ sb_1__8_.mux_bottom_track_25.out VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__284
+ VGND VGND VPWR VPWR net284 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__284/LO
+ sky130_fd_sc_hd__conb_1
X_272_ net62 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input76_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__A sb_1__8_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output232_A net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_1.mux_l2_in_0_ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput214 net214 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
Xoutput203 net203 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_2.mux_l4_in_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_0__S sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net278 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.out sky130_fd_sc_hd__buf_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_36.mux_l1_in_1_ net71 net83 sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__S cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__266__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_324_ net24 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk cby_1__8_.ccff_tail net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_2__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_29.mux_l1_in_2_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net74 sb_1__8_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ sb_1__8_.mem_bottom_track_25.ccff_tail net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_27.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_5.mux_l1_in_1__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_3_ net264 sb_1__8_.mux_bottom_track_45.out cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.out sky130_fd_sc_hd__buf_4
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input39_A chanx_right_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_1.mux_l1_in_1_ net222 net219 sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_31.mux_l1_in_0__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_7.mux_l2_in_3__351 VGND VGND VPWR VPWR net351 sb_1__8_.mux_left_track_7.mux_l2_in_3__351/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_1.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
X_307_ net8 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__370 VGND VGND VPWR VPWR net370 cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__370/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2_ net14 cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.mux_l3_in_1_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_7.mux_l2_in_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk sb_1__8_.mem_right_track_44.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__363 VGND VGND VPWR VPWR net363
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__363/LO sky130_fd_sc_hd__conb_1
XFILLER_88_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_2.mux_l2_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net304 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3_ net249 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_37.mux_l1_in_0_ net33 net44 sb_1__8_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_3__266 VGND VGND VPWR VPWR net266 cby_1__8_.mux_right_ipin_9.mux_l2_in_3__266/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_23.mux_l1_in_0__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_49.mux_l2_in_0_ net336 sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_49.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput114 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput103 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_2_ net86 cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3_ net38 net7 cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_0.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_left_track_7.mux_l1_in_1_ net70 net82 sb_1__8_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_51.mux_l2_in_0_ net338 sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_51.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__274__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_7.mux_l4_in_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__A1 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_3_ net256 net54 cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_3.mux_l2_in_2__A0 net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_3__S sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out net5
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_9.mux_l1_in_1__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__S cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__269__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2_ net30 net41 cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_94_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_29.mux_l2_in_0_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_3_ sb_1__8_.mux_bottom_track_29.out net69 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_0__S sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_85_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_head net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_340_ sb_1__8_.mux_bottom_track_27.out VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_271_ sb_1__8_.mux_left_track_45.out VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__287
+ VGND VGND VPWR VPWR net287 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__287/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_7.mux_l3_in_1_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input69_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3_ net364 net58 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_6__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output225_A net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2__A1 net35 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput215 net215 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
Xoutput204 net204 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput226 net226 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_36.mux_l1_in_0_ net105 net111 sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_19_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_323_ sb_1__8_.mux_right_track_0.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XANTENNA__282__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_13.mux_l4_in_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_29.mux_l1_in_1_ net66 net78 sb_1__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__301
+ VGND VGND VPWR VPWR net301 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__301/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_2__A0 sb_1__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_0.mux_l1_in_0_ net111 net108 sb_1__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_17.mux_l2_in_1__319 VGND VGND VPWR VPWR net319 sb_1__8_.mux_bottom_track_17.mux_l2_in_1__319/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__8_.mux_left_track_5.mux_l1_in_1__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_2_ net90 sb_1__8_.mux_bottom_track_27.out cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4_ net35 net4 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_1.mux_l1_in_0_ net224 net51 sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__277__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_31.mux_l1_in_0__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_306_ net7 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.mux_l3_in_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk sb_1__8_.mem_right_track_36.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__273
+ VGND VGND VPWR VPWR net273 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__273/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_13.mux_l3_in_1_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2__A0 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_34_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input51_A chanx_right_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_53.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_60_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_3__S sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput104 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__clkbuf_2
Xinput115 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net115
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_1_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_29_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_0.mux_l2_in_2__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l2_in_2__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_left_track_7.mux_l1_in_0_ net59 net46 sb_1__8_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input99_A reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__290__A sb_1__8_.mux_left_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_0__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4__A0 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_17.mux_l2_in_0__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk sb_1__8_.mem_bottom_track_7.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk sb_1__8_.mem_bottom_track_13.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_2_ net74 sb_1__8_.mux_bottom_track_39.out cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_3.mux_l2_in_2__A1 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_3__254 VGND VGND VPWR VPWR net254 cby_1__8_.mux_right_ipin_11.mux_l2_in_3__254/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_58_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_46_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mux_bottom_track_9.mux_l1_in_1__A1 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__285__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_49.mux_l1_in_0_ net222 net49 sb_1__8_.mem_bottom_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1_ net10 cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_39_prog_clk
+ sb_1__8_.mem_bottom_track_45.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_45.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_2_ sb_1__8_.mux_bottom_track_17.out net76 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_51.mux_l1_in_0_ net223 net50 sb_1__8_.mem_bottom_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_270_ net60 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_7.mux_l3_in_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2_ net27 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output218_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_58_prog_clk cby_1__8_.mem_right_ipin_1.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput216 net216 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput205 net205 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput227 net227 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_87_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_59_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2_ net48 net17 cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_322_ sb_1__8_.mux_right_track_2.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input81_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_29.mux_l1_in_0_ net44 net39 sb_1__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__285
+ VGND VGND VPWR VPWR net285 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__285/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_1_ net70 cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3_ net41 net10 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_0.mux_l2_in_3__352 VGND VGND VPWR VPWR net352 sb_1__8_.mux_right_track_0.mux_l2_in_3__352/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk sb_1__8_.mem_left_track_21.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__293__A sb_1__8_.mux_left_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_305_ sb_1__8_.mux_right_track_36.out VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net314 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net118 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3__A0 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_13.mux_l3_in_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_0__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A chanx_right_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__288__A sb_1__8_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk sb_1__8_.mem_left_track_53.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mux_right_ipin_7.mux_l1_in_2_ sb_1__8_.mux_bottom_track_15.out net77 cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_0__A0 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput105 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l2_in_2__A1 sb_1__8_.mux_bottom_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2__A0 net28 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_0__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4__A1 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_4.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l2_in_3__A1 sb_1__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_1__8_.mem_bottom_track_13.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_1_ net64 cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_46_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_88_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk
+ sb_1__8_.mem_bottom_track_43.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_45.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_2__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__A1 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__297
+ VGND VGND VPWR VPWR net297 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__297/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__296__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__276
+ VGND VGND VPWR VPWR net276 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__276/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_13.mux_l1_in_2_ sb_1__8_.mux_bottom_track_27.out net70 cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1__A0 sb_1__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput217 net217 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
Xoutput206 net206 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput228 net228 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__368 VGND VGND VPWR VPWR net368 cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__368/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk
+ sb_1__8_.mem_bottom_track_19.mem_out\[1\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_19.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_input109_A right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ sb_1__8_.mux_right_track_4.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input74_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_19.mux_l3_in_0_ sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_19.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_output230_A net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_25.mux_l1_in_1__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_45_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_45.mux_l1_in_0__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_1__8_.mem_left_track_21.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_304_ net5 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3__A1 net11 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_7.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_0__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_19.mux_l2_in_1_ net320 net3 sb_1__8_.mem_bottom_track_19.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_20.mux_l1_in_3_ net356 net25 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input37_A chanx_right_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_86_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk sb_1__8_.mem_left_track_45.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_1__S sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_7.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__306
+ VGND VGND VPWR VPWR net306 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__306/LO
+ sky130_fd_sc_hd__conb_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput106 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__248 VGND VGND VPWR VPWR net248 cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__248/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__299__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_1__8_.mem_bottom_track_11.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_11.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_20.mux_l3_in_0_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_2__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2__A0 sb_1__8_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_13.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xoutput207 net207 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput229 net229 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_53.mux_l1_in_0__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_3.mux_l2_in_3_ net346 net233 sb_1__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_1__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l2_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk
+ sb_1__8_.mem_bottom_track_19.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_19.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_320_ sb_1__8_.mux_right_track_6.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__A0 sb_1__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input67_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output223_A net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_20.mux_l2_in_1_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_left_track_45.mux_l1_in_0__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xsb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__8_.mem_right_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__269
+ VGND VGND VPWR VPWR net269 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__269/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_2.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk sb_1__8_.mem_left_track_13.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
X_303_ net4 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_0__A0 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_5.mux_l2_in_3__A1 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_19.mux_l2_in_0_ net7 sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_19.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_20.mux_l1_in_2_ net11 net87 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_3.mux_l4_in_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_13.mux_l1_in_3_ net343 net229 sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_7.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_21.mux_l2_in_0_ sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput107 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_29.mux_l1_in_0__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_1__S sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net295 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_3.mux_l3_in_1_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l1_in_2__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input97_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_21.mux_l1_in_1_ net321 net5 sb_1__8_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net267 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_6.mux_l2_in_3_ net362 net29 sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_13.mux_l3_in_0_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_0.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_13.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput208 net208 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__8_.mux_left_track_53.mux_l1_in_0__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_3.mux_l2_in_2_ net230 net227 sb_1__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net300 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__mux2_4
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk
+ sb_1__8_.mem_bottom_track_17.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_19.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_20.mux_l2_in_0_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_44.mux_l2_in_1__360 VGND VGND VPWR VPWR net360 sb_1__8_.mux_right_track_44.mux_l2_in_1__360/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_13.mux_l2_in_1_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out
+ net23 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk sb_1__8_.mem_right_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l2_in_3__A1 sb_1__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input114_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ net236 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfrtp_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mux_bottom_track_19.mux_l2_in_1__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__271
+ VGND VGND VPWR VPWR net271 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__271/LO
+ sky130_fd_sc_hd__conb_1
X_302_ net32 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xsb_1__8_.mux_right_track_6.mux_l4_in_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_0__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_1__8_.mem_bottom_track_31.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_2__S sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_3__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_20.mux_l1_in_1_ net69 net81 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_3__264 VGND VGND VPWR VPWR net264 cby_1__8_.mux_right_ipin_7.mux_l2_in_3__264/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_3__A1 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_13.mux_l1_in_2_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net86 sb_1__8_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__S cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_49.mux_l2_in_0__336 VGND VGND VPWR VPWR net336 sb_1__8_.mux_bottom_track_49.mux_l2_in_0__336/LO
+ sky130_fd_sc_hd__conb_1
Xinput108 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND
+ VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_6.mux_l3_in_1_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_29.mux_l1_in_0__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_right_track_44.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__A0 sb_1__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input42_A chanx_right_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk cby_1__8_.mem_right_ipin_3.ccff_tail
+ net237 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_19.mux_l1_in_0_ net219 net37 sb_1__8_.mem_bottom_track_19.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_38_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_6.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_3.mux_l3_in_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput90 chany_bottom_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
Xsb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_41_prog_clk
+ sb_1__8_.mem_bottom_track_37.mem_out\[1\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_37.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_21.mux_l1_in_0_ net220 net35 sb_1__8_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_0__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3__A0 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_33.mux_l2_in_0_ net328 sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_33.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_11.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_6.mux_l2_in_2_ net16 net74 sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1__A0 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_89_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput209 net209 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_3.mux_l2_in_1_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net90 sb_1__8_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_6.mux_l1_in_3_ net66 net78 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_45.mux_l1_in_0__A0 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_13.mux_l2_in_0_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__S cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_1__S sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input107_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_301_ sb_1__8_.mux_right_track_44.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input72_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_6.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ sb_1__8_.mem_bottom_track_29.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_31.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_45.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_2__S sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__302__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_bottom_track_37.mux_l1_in_0__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_right_track_52.mux_l1_in_0__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_20.mux_l1_in_0_ net103 net109 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net284 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__267
+ VGND VGND VPWR VPWR net267 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__267/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_13.mux_l1_in_1_ net68 net80 sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_2__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2__A0 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput109 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND
+ VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_1__8_.mux_right_track_44.mux_l3_in_0_ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_6.mux_l3_in_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_44.mux_l1_in_0__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_79_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input35_A chanx_right_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3_ net240 net60 cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_7.mux_l3_in_0_ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_3.mux_l1_in_0__A0 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_right_track_6.mux_l2_in_2__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__281
+ VGND VGND VPWR VPWR net281 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__281/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput80 chany_bottom_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
Xinput91 chany_bottom_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk
+ sb_1__8_.mem_bottom_track_37.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_37.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net285 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_44.mux_l2_in_1_ net360 sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_right_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_6.mux_l2_in_1_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__310__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_1.mux_l1_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_3_ net260 net53 cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_7.mux_l2_in_1_ net339 sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l2_in_3__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_3.mux_l2_in_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_1.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__A1 net44 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3_ net245 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net282 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__mux2_4
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_44.mux_l1_in_2_ net7 net90 sb_1__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_bottom_track_33.mux_l1_in_0_ net26 net56 sb_1__8_.mem_bottom_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_6.mux_l1_in_2_ net106 net104 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_3__A0 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk sb_1__8_.mem_left_track_13.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_45.mux_l2_in_0_ net334 sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_45.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_15.mux_l2_in_1__318 VGND VGND VPWR VPWR net318 sb_1__8_.mux_bottom_track_15.mux_l2_in_1__318/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__279
+ VGND VGND VPWR VPWR net279 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__279/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__8_.mux_bottom_track_7.mux_l1_in_2_ net16 net19 sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__311
+ VGND VGND VPWR VPWR net311 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__311/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_300_ net30 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_11.mux_l1_in_0__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_3.mux_l1_in_1_ net72 net84 sb_1__8_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input65_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net114 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output221_A net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_3.mux_l4_in_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk sb_1__8_.mem_left_track_45.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 ccff_head_1 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_right_track_52.mux_l1_in_0__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4_ net34 net32 cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_sb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_left_track_11.mux_l2_in_2__A0 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_13.mux_l1_in_0_ net56 net42 sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_4.mem_out\[2\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_80_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_3_ net265 net52 cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_37.mux_l3_in_0_ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput190 net190 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2_ net29 net37 cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_3.mux_l3_in_1_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_bottom_track_3.mux_l1_in_0__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__308__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 chany_bottom_in[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
Xinput81 chany_bottom_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput92 chany_bottom_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ sb_1__8_.mem_bottom_track_35.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_37.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3_ net250 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_4_ sb_1__8_.mux_bottom_track_41.out net92 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_44.mux_l2_in_0_ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_6.mux_l2_in_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_1.mux_l1_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_37.mux_l2_in_1_ net347 sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_2_ net85 sb_1__8_.mux_bottom_track_37.out cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_7.mux_l2_in_0_ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input95_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_8.mux_l4_in_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk cby_1__8_.mem_right_ipin_10.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_3_ net257 net52 cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_0__S sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_1.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.out sky130_fd_sc_hd__buf_4
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__A0 sb_1__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1__A0 sb_1__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2_ net26 cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_44.mux_l1_in_1_ net72 net84 sb_1__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_6.mux_l1_in_1_ net102 net100 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_3__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_37.mux_l1_in_2_ net232 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__8_.mem_left_track_37.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk sb_1__8_.mem_left_track_13.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_7.mux_l1_in_1_ net222 net219 sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA__316__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A ccff_head_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_8.mux_l3_in_1_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3_ net365 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net311 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__mux2_4
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_7.mux_l2_in_1__339 VGND VGND VPWR VPWR net339 sb_1__8_.mux_bottom_track_7.mux_l2_in_1__339/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_50_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_11.mux_l1_in_0__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_3.mux_l1_in_0_ net62 net48 sb_1__8_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_4_ sb_1__8_.mux_bottom_track_41.out net92 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A chanx_right_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l2_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_5.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_359_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk sb_1__8_.mem_left_track_37.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 ccff_head_2 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3_ sb_1__8_.mux_left_track_29.out net9
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_19_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_14.mux_l4_in_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_left_track_11.mux_l2_in_2__A1 net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input112_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__A0 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_45.mux_l1_in_0_ net220 net40 sb_1__8_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_2_ net86 cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__310
+ VGND VGND VPWR VPWR net310 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__310/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__246 VGND VGND VPWR VPWR net246 cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__246/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput191 net191 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput180 net180 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_1_ net6 cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_3.mux_l3_in_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_1__S sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_13.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew235 net238 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_3__S sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__324__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_14.mux_l3_in_1_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xinput71 chany_bottom_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput82 chany_bottom_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 net112 net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2_ net14 net35 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__270
+ VGND VGND VPWR VPWR net270 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__270/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mem_bottom_track_41.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input40_A chanx_right_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_3_ sb_1__8_.mux_bottom_track_29.out net69 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_16_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net303 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_59_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_37.mux_l2_in_0_ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__319__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_1_ net65 cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input88_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_2_ net86 cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net274 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_0__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_44.mux_l1_in_0_ net106 net100 sb_1__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_28.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_57_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_6.mux_l1_in_0_ net110 net108 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_11.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_left_track_37.mux_l1_in_1_ net63 net65 sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_3.mux_l1_in_2_ sb_1__8_.mux_bottom_track_19.out net75 cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_48_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_7.mux_l1_in_0_ net224 net46 sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_8.mux_l3_in_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2_ net26 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__300
+ VGND VGND VPWR VPWR net300 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__300/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_3_ sb_1__8_.mux_bottom_track_29.out net69 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_5.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_358_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mux_bottom_track_5.mux_l1_in_1__A0 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ net51 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__327__A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input105_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2__A0 net27 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input70_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_4.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l2_in_3__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_1_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3_ sb_1__8_.mux_left_track_29.out
+ net9 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2__A1 net39 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_3__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput170 net170 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew236 net98 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_12
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l1_in_1__A0 sb_1__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_14.mux_l3_in_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 chany_bottom_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xinput83 chany_bottom_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1_ net4 cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_35.mux_l2_in_0__329 VGND VGND VPWR VPWR net329 sb_1__8_.mux_bottom_track_35.mux_l2_in_0__329/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input33_A chanx_right_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_2_ sb_1__8_.mux_bottom_track_17.out net76 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_15.mux_l3_in_0_ sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_15.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_10.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__335__A sb_1__8_.mux_bottom_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_3__251 VGND VGND VPWR VPWR net251 cby_1__8_.mux_right_ipin_0.mux_l2_in_3__251/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_1_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2_ net41 net10 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3__A0 net38 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_15.mux_l2_in_1_ net318 net31 sb_1__8_.mem_bottom_track_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk sb_1__8_.mem_right_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__289
+ VGND VGND VPWR VPWR net289 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__289/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_1__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_37.mux_l1_in_0_ net77 net38 sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_3.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_1.mux_l2_in_2__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_13.mux_l2_in_0__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk
+ sb_1__8_.mem_bottom_track_23.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_23.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_2_ sb_1__8_.mux_bottom_track_17.out net76 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_1__8_.mem_left_track_5.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_65_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_357_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_bottom_track_5.mux_l1_in_1__A1 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_288_ sb_1__8_.mux_left_track_11.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net293 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__mux2_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_3__262 VGND VGND VPWR VPWR net262 cby_1__8_.mux_right_ipin_5.mux_l2_in_3__262/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input63_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_2.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_3__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput160 net160 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput171 net171 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew237 net98 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_12
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_46_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xinput73 chany_bottom_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xinput84 chany_bottom_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__A0 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2__A0 net41 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__8_.mem_bottom_track_5.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_2__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__366 VGND VGND VPWR VPWR net366
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__366/LO sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__8_.mux_right_track_10.mux_l2_in_2__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_2__S sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__242 VGND VGND VPWR VPWR net242 cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__242/LO
+ sky130_fd_sc_hd__conb_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_0__S sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_10.ccff_head
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_3__259 VGND VGND VPWR VPWR net259 cby_1__8_.mux_right_ipin_2.mux_l2_in_3__259/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net292 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net301 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_15.mux_l2_in_0_ net9 sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_15.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk sb_1__8_.mem_right_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_45_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input93_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_2.mux_l1_in_0__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_3.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2__A0 net26 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ sb_1__8_.mem_bottom_track_21.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_23.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk sb_1__8_.mem_left_track_37.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_5.mux_l1_in_0__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_29_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk sb_1__8_.mem_left_track_3.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_356_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_287_ sb_1__8_.mux_left_track_13.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input56_A chanx_right_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__296
+ VGND VGND VPWR VPWR net296 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__296/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_339_ sb_1__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out
+ net19 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_47.mux_l2_in_0__335 VGND VGND VPWR VPWR net335 sb_1__8_.mux_bottom_track_47.mux_l2_in_0__335/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_2.mux_l2_in_3_ net355 net32 sb_1__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_3__S sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput161 net161 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input110_A right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_0.mux_l2_in_1__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_1__8_.mem_bottom_track_29.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__264__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_12.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew238 net98 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_12
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_46_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xinput63 chany_bottom_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput85 chany_bottom_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput74 chany_bottom_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_21.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_3.mux_l2_in_1__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_5.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_9.mux_l1_in_0__A0 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_2.mux_l4_in_0_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sb_1__8_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_75_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_7.mux_l1_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l2_in_3__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input86_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__272__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_3__257 VGND VGND VPWR VPWR net257 cby_1__8_.mux_right_ipin_14.mux_l2_in_3__257/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk sb_1__8_.mem_left_track_37.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_1__S sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_5.mux_l1_in_0__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_2.mux_l3_in_1_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__S cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_355_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_286_ net48 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_15.mux_l1_in_0_ net225 net39 sb_1__8_.mem_bottom_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_17.mux_l1_in_0__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_27.mux_l2_in_0_ sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_27.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input49_A chanx_right_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net275 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__mux2_4
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_338_ sb_1__8_.mux_bottom_track_31.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_left_track_21.mux_l1_in_3_ net344 net230 sb_1__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_269_ net59 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XANTENNA_load_slew239_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out
+ net22 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_2.mux_l2_in_2_ net18 net64 sb_1__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput151 net151 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_0.mux_l2_in_1__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input103_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l2_in_1__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_27.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__280__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3__A0 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xload_slew239 net98 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_12
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_46_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xinput64 chany_bottom_in[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__D cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xinput86 chany_bottom_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xinput75 chany_bottom_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__313
+ VGND VGND VPWR VPWR net313 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__313/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_left_track_3.mux_l2_in_1__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_27.mux_l1_in_1_ net324 net30 sb_1__8_.mem_bottom_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_3.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_bottom_track_9.mux_l1_in_0__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net290 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_41.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk
+ sb_1__8_.mem_bottom_track_41.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_41.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_3__A1 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_21.mux_l3_in_0_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_bottom_track_7.mux_l1_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net310 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_1__S sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input79_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_25.mux_l1_in_0__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_13.mux_l2_in_1__317 VGND VGND VPWR VPWR net317 sb_1__8_.mux_bottom_track_13.mux_l2_in_1__317/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_21.mux_l2_in_1_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_29.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_2.mux_l3_in_0_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_5.mux_l2_in_1__337 VGND VGND VPWR VPWR net337 sb_1__8_.mux_bottom_track_5.mux_l2_in_1__337/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_51.mux_l2_in_0__338 VGND VGND VPWR VPWR net338 sb_1__8_.mux_bottom_track_51.mux_l2_in_0__338/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_354_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__283__A sb_1__8_.mux_left_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ net47 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_3.mux_l3_in_0_ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l1_in_2__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2__A0 sb_1__8_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_bottom_track_17.mux_l1_in_0__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__308
+ VGND VGND VPWR VPWR net308 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__308/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__278__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_1__8_.mux_bottom_track_33.out VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_21.mux_l1_in_2_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net85 sb_1__8_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_268_ net58 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_2.mux_l2_in_1_ net76 net106 sb_1__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_37_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__A0 sb_1__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput141 net141 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__244 VGND VGND VPWR VPWR net244 cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__244/LO
+ sky130_fd_sc_hd__conb_1
Xoutput174 net174 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput196 net196 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.out sky130_fd_sc_hd__clkbuf_2
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_3.mux_l2_in_1_ net326 sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input61_A chanx_right_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3__A1 net10 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__304
+ VGND VGND VPWR VPWR net304 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__304/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_46_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xinput76 chany_bottom_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput65 chany_bottom_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput87 chany_bottom_in[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput98 prog_reset VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_0.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_27.mux_l1_in_0_ net223 net60 sb_1__8_.mem_bottom_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__8_.mux_right_track_4.mux_l1_in_1__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_39.mux_l2_in_0_ net331 sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_39.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3_ net367 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__291__A sb_1__8_.mux_left_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l2_in_3__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_15.mux_l2_in_1__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_41.mux_l2_in_0_ net332 sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_41.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_41.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk
+ sb_1__8_.mem_bottom_track_39.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_41.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_3.mux_l1_in_2_ net18 net22 sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3_ net241 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_bottom_track_33.mux_l1_in_0__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__286__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0__A0 sb_1__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_29.mux_l2_in_0__325 VGND VGND VPWR VPWR net325 sb_1__8_.mux_bottom_track_29.mux_l2_in_0__325/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4_ sb_1__8_.mux_left_track_45.out net30
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_1__8_.mem_bottom_track_15.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output228_A net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_25.mux_l1_in_0__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_42_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_21.mux_l2_in_0_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out net5
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_3_ net261 net54 cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_5__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_2.mux_l2_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk
+ sb_1__8_.mem_bottom_track_47.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_47.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_353_ sb_1__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
X_284_ net46 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input91_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__299
+ VGND VGND VPWR VPWR net299 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__299/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_5.mux_l2_in_2__A0 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_3.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3_ net246 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__294__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ sb_1__8_.mux_bottom_track_35.out VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_left_track_21.mux_l1_in_1_ net67 net79 sb_1__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_4_ sb_1__8_.mux_bottom_track_45.out net90 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
X_267_ sb_1__8_.mux_left_track_53.out VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_2.mux_l2_in_0_ net103 sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__A1 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput120 net120 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_right_track_52.mux_l3_in_0_ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xoutput197 net197 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_3.mux_l2_in_0_ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input54_A chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l4_in_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA__289__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_47_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_3_ net253 net54 cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
X_319_ net21 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput77 chany_bottom_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
Xinput66 chany_bottom_in[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xinput88 chany_bottom_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_4
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xinput99 reset VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.out sky130_fd_sc_hd__buf_4
XFILLER_69_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_41.mux_l1_in_0__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_4.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2_ net14 cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l1_in_1__A0 sb_1__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_3_ net266 sb_1__8_.mux_bottom_track_49.out cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__A1 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_52.mux_l2_in_1_ net361 net5 sb_1__8_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_1__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_bottom_track_3.mux_l1_in_1_ net223 net220 sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_45.mux_l2_in_1__348 VGND VGND VPWR VPWR net348 sb_1__8_.mux_left_track_45.mux_l2_in_1__348/LO
+ sky130_fd_sc_hd__conb_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_4.mux_l3_in_1_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_33.mux_l1_in_0__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_4_ sb_1__8_.mux_bottom_track_45.out net90 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ net236 VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_39.mux_l1_in_0_ net225 net57 sb_1__8_.mem_bottom_track_39.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3_ net38 net7 cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_6.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_10.mux_l4_in_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_1__8_.mem_bottom_track_15.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3__A0 net38 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_41.mux_l1_in_0_ net218 net61 sb_1__8_.mem_bottom_track_41.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_76_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net271 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_11_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_2_ net74 cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mux_right_track_2.mux_l2_in_2__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l2_in_2__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_9.mux_l4_in_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_85_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk
+ sb_1__8_.mem_bottom_track_45.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_47.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_352_ sb_1__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4__A0 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_19.mux_l2_in_0__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_283_ sb_1__8_.mux_left_track_21.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input84_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_3_ net258 sb_1__8_.mux_bottom_track_43.out
+ cby_1__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_5.mux_l2_in_2__A1 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_57_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_10.mux_l3_in_1_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2_ net28 net39 cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_51_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_10.mux_l2_in_3_ net353 net28 sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_3__260 VGND VGND VPWR VPWR net260 cby_1__8_.mux_right_ipin_3.mux_l2_in_3__260/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_335_ sb_1__8_.mux_bottom_track_37.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_left_track_21.mux_l1_in_0_ net55 net41 sb_1__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_3_ sb_1__8_.mux_bottom_track_33.out net67 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_266_ net56 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_2__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_60_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_9.mux_l3_in_1_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3_ net366 net56 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xoutput132 net132 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net312 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__mux2_4
Xoutput165 net165 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput198 net198 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_45.mux_l3_in_0_ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input47_A chanx_right_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_47_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_2__S sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_2_ net74 cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
X_318_ sb_1__8_.mux_right_track_10.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput78 chany_bottom_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput67 chany_bottom_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
Xinput89 chany_bottom_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XANTENNA_load_slew237_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_15.mux_l4_in_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.ccff_tail VGND
+ VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__371 VGND VGND VPWR VPWR net371 cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__371/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_33.mux_l2_in_0__328 VGND VGND VPWR VPWR net328 sb_1__8_.mux_bottom_track_33.mux_l2_in_0__328/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input101_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_9.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_2.mux_l1_in_0_ net100 net109 sb_1__8_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__364 VGND VGND VPWR VPWR net364
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__364/LO sky130_fd_sc_hd__conb_1
XFILLER_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_2_ net88 sb_1__8_.mux_bottom_track_31.out cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__240 VGND VGND VPWR VPWR net240 cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__240/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_47_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4_ net62 net31 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_52.mux_l2_in_0_ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_right_track_10.mux_l4_in_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_3.mux_l1_in_0_ net225 net48 sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_45.mux_l2_in_1_ net348 net233 sb_1__8_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l3_in_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_3_ sb_1__8_.mux_bottom_track_33.out net67 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_15.mux_l3_in_1_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_81_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk sb_1__8_.mem_bottom_track_13.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_70_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_1__8_.mem_left_track_29.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_10.mux_l3_in_1_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_52.mux_l1_in_1_ net91 net73 sb_1__8_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_6.mux_l2_in_3__362 VGND VGND VPWR VPWR net362 sb_1__8_.mux_right_track_6.mux_l2_in_3__362/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_1_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_left_track_5.mux_l2_in_3__349 VGND VGND VPWR VPWR net349 sb_1__8_.mux_left_track_5.mux_l2_in_3__349/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_2__A0 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_351_ sb_1__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4__A1 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_282_ net43 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_2_ net91 sb_1__8_.mux_bottom_track_31.out cby_1__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_input77_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output233_A net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l2_in_3__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail net97 VGND
+ VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_10.mux_l3_in_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__288
+ VGND VGND VPWR VPWR net288 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__288/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1_ net8 cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xsb_1__8_.mux_right_track_10.mux_l2_in_2_ net13 net85 sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net115 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_2__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ sb_1__8_.mux_bottom_track_39.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_2_ sb_1__8_.mux_bottom_track_21.out net73 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_265_ net55 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_11.mux_l3_in_0_ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_2__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_9.mux_l3_in_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2_ net25 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput133 net133 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__A1 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput177 net177 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__A0 sb_1__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_47_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_317_ sb_1__8_.mux_right_track_12.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_1_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
XFILLER_52_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput68 chany_bottom_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xinput79 chany_bottom_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net1
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2_ net46 net15 cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_10.mux_l1_in_3_ net67 net79 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_11.mux_l2_in_1_ net316 net10 sb_1__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_bottom_track_27.mux_l1_in_1__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_2__S sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2__A0 sb_1__8_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_1_ net68 cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__283
+ VGND VGND VPWR VPWR net283 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__283/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3_ net39 net8 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net117 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mux_right_ipin_11.mux_l2_in_1__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_0__S sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_45.mux_l2_in_0_ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_2_ sb_1__8_.mux_bottom_track_21.out net73 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l3_in_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_29.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_9.mux_l1_in_2_ sb_1__8_.mux_bottom_track_19.out net75 cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2__A0 net3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_10.mux_l3_in_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_52.mux_l1_in_0_ net107 net101 sb_1__8_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_76_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_3__255 VGND VGND VPWR VPWR net255 cby_1__8_.mux_right_ipin_12.mux_l2_in_3__255/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_71_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_45.mux_l1_in_1_ net227 net64 sb_1__8_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ sb_1__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_2__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_281_ net42 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_1_ net68 cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_2.ccff_tail
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net307 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_10.mux_l2_in_1_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_2__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net273 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ sb_1__8_.mux_bottom_track_41.out VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_264_ net44 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_45.mux_l2_in_0__334 VGND VGND VPWR VPWR net334 sb_1__8_.mux_bottom_track_45.mux_l2_in_0__334/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1__A0 sb_1__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_3__S sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput134 net134 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
XFILLER_87_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__278
+ VGND VGND VPWR VPWR net278 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__278/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_15.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mux_right_ipin_11.mux_l1_in_2__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail net97 VGND
+ VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
X_316_ net18 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_27.mux_l1_in_1__324 VGND VGND VPWR VPWR net324 sb_1__8_.mux_bottom_track_27.mux_l1_in_1__324/LO
+ sky130_fd_sc_hd__conb_1
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_4
Xsb_1__8_.mux_bottom_track_37.mux_l2_in_1__330 VGND VGND VPWR VPWR net330 sb_1__8_.mux_bottom_track_37.mux_l2_in_1__330/LO
+ sky130_fd_sc_hd__conb_1
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
Xinput69 chany_bottom_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net294 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__mux2_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_10.mux_l1_in_2_ net107 net105 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__S cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_11.mux_l2_in_0_ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_1__8_.mem_bottom_track_33.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_33.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_27_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input52_A chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_0__S sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_1.mux_l1_in_1__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_0__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_left_track_7.mux_l2_in_3__A1 net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_11.mux_l1_in_1_ net12 net221 sb_1__8_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk cby_1__8_.mem_right_ipin_5.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_80_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk sb_1__8_.mem_left_track_21.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_9.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2__A1 net34 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_45.mux_l1_in_0_ net76 net37 sb_1__8_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_2__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__290
+ VGND VGND VPWR VPWR net290 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__290/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_60_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ net41 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output219_A net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_45.mux_l2_in_1__A1 net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_10.mux_l2_in_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_2__S sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ sb_1__8_.mux_bottom_track_43.out VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input82_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_1__8_.mem_right_track_0.mem_out\[2\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput124 net124 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_3__S sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput135 net135 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
XANTENNA__303__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput157 net157 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
XFILLER_87_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput179 net179 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_5.mux_l2_in_3_ net349 net234 sb_1__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_56_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_315_ net17 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_10.mux_l1_in_1_ net103 net101 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_0__A0 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_8.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_43_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ sb_1__8_.mem_bottom_track_31.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_33.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input45_A chanx_right_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out
+ net21 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_load_slew235_A net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_2__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_1.mux_l1_in_1__A1 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l2_in_3__A1 sb_1__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_0__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__249 VGND VGND VPWR VPWR net249 cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__249/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l1_in_1__A0 sb_1__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_39.mux_l1_in_0__A0 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_11.mux_l1_in_0_ net218 net42 sb_1__8_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_5.mux_l4_in_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0__A0 sb_1__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_9.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_23.mux_l2_in_0_ sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_23.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net296 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mux_left_track_53.mux_l2_in_1__A1 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mem_bottom_track_39.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk
+ sb_1__8_.mem_bottom_track_39.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_39.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_2__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_11.mux_l2_in_1__316 VGND VGND VPWR VPWR net316 sb_1__8_.mux_bottom_track_11.mux_l2_in_1__316/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA__306__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_5.mux_l3_in_1_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_1.mem_out\[2\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_23.mux_l1_in_1_ net322 net4 sb_1__8_.mem_bottom_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_331_ sb_1__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net291 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_44.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input75_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output231_A net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_1__8_.mem_right_track_0.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput125 net125 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_36_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_5.mux_l2_in_2_ net231 net228 sb_1__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_86_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_314_ net16 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_2__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_10.mux_l1_in_0_ net111 net109 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__sdfrtp_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__314__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_0__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net276 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__mux2_4
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input38_A chanx_right_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_1.mux_l1_in_0__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out
+ net24 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_47.mux_l1_in_0__A0 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_6.mem_out\[2\]
+ net239 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_21.mux_l1_in_3__344 VGND VGND VPWR VPWR net344 sb_1__8_.mux_left_track_21.mux_l1_in_3__344/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.out sky130_fd_sc_hd__buf_4
XFILLER_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__293
+ VGND VGND VPWR VPWR net293 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__293/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__302
+ VGND VGND VPWR VPWR net302 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__302/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_39.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk
+ sb_1__8_.mem_bottom_track_37.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_39.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_19.mux_l2_in_1__320 VGND VGND VPWR VPWR net320 sb_1__8_.mux_bottom_track_19.mux_l2_in_1__320/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_79_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2__A0 sb_1__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_1__S sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_3.mux_l2_in_3__346 VGND VGND VPWR VPWR net346 sb_1__8_.mux_left_track_3.mux_l2_in_3__346/LO
+ sky130_fd_sc_hd__conb_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_3.mux_l2_in_1__326 VGND VGND VPWR VPWR net326 sb_1__8_.mux_bottom_track_3.mux_l2_in_1__326/LO
+ sky130_fd_sc_hd__conb_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_5.mux_l3_in_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_1.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_71_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_5.mux_l1_in_0__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_4__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_23.mux_l1_in_0_ net221 net34 sb_1__8_.mem_bottom_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_12.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk
+ sb_1__8_.mem_bottom_track_51.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_51.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
X_330_ sb_1__8_.mux_bottom_track_47.out VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_35.mux_l2_in_0_ net329 sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_35.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_44.mux_l1_in_2__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input68_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output224_A net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_27_prog_clk sb_1__8_.mem_right_track_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_37.mux_l2_in_1__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput137 net137 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__8_.mux_bottom_track_3.mux_l1_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3_ net369 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_5.mux_l2_in_1_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net89 sb_1__8_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l2_in_3__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_313_ sb_1__8_.mux_right_track_20.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XANTENNA_sb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk sb_1__8_.mem_left_track_7.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__A1 sb_1__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_left_track_1.mux_l1_in_0__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_2__S sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_3_ net251 sb_1__8_.mux_bottom_track_49.out cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4_ net34 net32 cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__325__A net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_6.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_3__265 VGND VGND VPWR VPWR net265 cby_1__8_.mux_right_ipin_8.mux_l2_in_3__265/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net305 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__mux2_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_13.mux_l1_in_0__A0 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input50_A chanx_right_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2__A0 sb_1__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3_ net368 net44 cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk cby_1__8_.mem_right_ipin_15.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR cby_1__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input98_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_20.mux_l1_in_3__356 VGND VGND VPWR VPWR net356 sb_1__8_.mux_right_track_20.mux_l1_in_3__356/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_4_ sb_1__8_.mux_bottom_track_37.out net65 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mux_right_ipin_1.mux_l2_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2__A1 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3_ net242 net58 cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_9.mux_l3_in_0_ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_0.mux_l4_in_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_1__8_.mem_left_track_1.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_5.mux_l1_in_0__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_12.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__333__A sb_1__8_.mux_bottom_track_41.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk
+ sb_1__8_.mem_bottom_track_49.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_51.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net309 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk net2
+ net239 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net277 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_3_ net262 net24 cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput116 net116 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__8_.mux_right_track_52.mux_l2_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput138 net138 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_9.mux_l2_in_1_ net340 sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_9.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_3.mux_l1_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_2__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2_ net26 cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_0.mux_l3_in_1_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_5.mux_l2_in_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input115_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_312_ net13 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input80_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net280 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__280
+ VGND VGND VPWR VPWR net280 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__280/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3_ net247 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk sb_1__8_.mem_left_track_7.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_21.mux_l1_in_0__A0 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_35.mux_l1_in_0_ net25 net55 sb_1__8_.mem_bottom_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_31.mux_l2_in_0__327 VGND VGND VPWR VPWR net327 sb_1__8_.mux_bottom_track_31.mux_l2_in_0__327/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__8_.mem_bottom_track_1.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_47.mux_l2_in_0_ net335 sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_47.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_3__A1 net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_9.mux_l1_in_2_ net13 net15 sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_2_ net88 cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3_ sb_1__8_.mux_left_track_29.out net9
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_sb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_5.mux_l1_in_1_ net71 net83 sb_1__8_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_6.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__8_.mux_right_ipin_1.mux_l1_in_2__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_55_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2__A0 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_13.mux_l1_in_0__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_5.mux_l4_in_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input43_A chanx_right_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_3_ net254 net52 cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4_ sb_1__8_.mux_left_track_45.out net30
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_bottom_track_43.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2_ net3 net34 cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk cby_1__8_.mem_right_ipin_15.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_3__253 VGND VGND VPWR VPWR net253 cby_1__8_.mux_right_ipin_10.mux_l2_in_3__253/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__282
+ VGND VGND VPWR VPWR net282 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__282/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_3_ sb_1__8_.mux_bottom_track_25.out net71 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_62_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_5.mux_l3_in_1_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2_ net27 net35 cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_1.mux_l2_in_3__341 VGND VGND VPWR VPWR net341 sb_1__8_.mux_left_track_1.mux_l2_in_3__341/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_81_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_1_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_1__8_.mem_bottom_track_51.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_0__S sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_11.mux_l4_in_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_bottom_track_11.mux_l2_in_1__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__292
+ VGND VGND VPWR VPWR net292 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__292/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_3.mux_l1_in_1__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_2_ net63 sb_1__8_.mux_bottom_track_41.out cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput139 net139 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_bottom_track_9.mux_l2_in_0_ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_0.mux_l3_in_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_21.mux_l1_in_3__A1 net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input108_A right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_0.mux_l2_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_311_ net12 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk sb_1__8_.mem_right_track_10.mem_out\[2\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input73_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ sb_1__8_.mem_bottom_track_25.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_25.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__312
+ VGND VGND VPWR VPWR net312 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__312/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_11.mux_l3_in_1_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2_ net14 cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk sb_1__8_.mem_left_track_7.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_21.mux_l1_in_0__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_39.mux_l2_in_0__331 VGND VGND VPWR VPWR net331 sb_1__8_.mux_bottom_track_39.mux_l2_in_0__331/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_8.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_9.mux_l1_in_1_ net223 net220 sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_42_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_1_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_left_track_5.mux_l1_in_0_ net60 net47 sb_1__8_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_4.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_2__A0 net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_2_ net86 sb_1__8_.mux_bottom_track_35.out cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_input36_A chanx_right_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_7.mux_l1_in_1__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3_ net38 net7 cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net287 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__mux2_4
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1_ net32 cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_47.mux_l1_in_0_ net221 net45 sb_1__8_.mem_bottom_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA__352__A sb_1__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_1__S sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk sb_1__8_.mem_bottom_track_7.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2__A1 net37 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1_ net4 cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_5.mux_l3_in_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2_ net43 net12 cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_11.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_31_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__275
+ VGND VGND VPWR VPWR net275 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__275/LO
+ sky130_fd_sc_hd__conb_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_3.mux_l1_in_1__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__367 VGND VGND VPWR VPWR net367 cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__367/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__A0 sb_1__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_1_ net92 cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_43.mux_l2_in_0__333 VGND VGND VPWR VPWR net333 sb_1__8_.mux_bottom_track_43.mux_l2_in_0__333/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_17_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput129 net129 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__250 VGND VGND VPWR VPWR net250 cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__250/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_310_ net11 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_1__8_.mem_right_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_53.mux_l3_in_0_ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input66_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ sb_1__8_.mem_bottom_track_23.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_25.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__270__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2__A0 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_25.mux_l1_in_1__323 VGND VGND VPWR VPWR net323 sb_1__8_.mux_bottom_track_25.mux_l1_in_1__323/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net298 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output222_A net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_11.mux_l3_in_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_5.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net313 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk sb_1__8_.mem_bottom_track_1.ccff_head
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_5.mux_l1_in_2_ sb_1__8_.mux_bottom_track_23.out net72 cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__S cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_9.mux_l1_in_0_ net225 net43 sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__265__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l2_in_2__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mem_bottom_track_39.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_bottom_track_15.mux_l2_in_0__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_53.mux_l2_in_1_ net350 net234 sb_1__8_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_2__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__305
+ VGND VGND VPWR VPWR net305 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__305/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_1_ net66 cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_7.mux_l1_in_1__A1 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__247 VGND VGND VPWR VPWR net247 cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__247/LO
+ sky130_fd_sc_hd__conb_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_14.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_sb_1__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__303
+ VGND VGND VPWR VPWR net303 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__303/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_right_track_12.mux_l1_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_11.mux_l1_in_2_ sb_1__8_.mux_bottom_track_23.out net72 cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__272
+ VGND VGND VPWR VPWR net272 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__272/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input96_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__273__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_2__S sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_12.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_17.mux_l3_in_0_ sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_17.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_26_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3__S cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_11.mux_l2_in_3_ net342 net234 sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__268__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput119 net119 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3__A0 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l1_in_4__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_1__8_.mem_right_track_10.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_10_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chanx_right_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail
+ net236 VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_17.mux_l2_in_1_ net319 net27 sb_1__8_.mem_bottom_track_17.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_1__8_.mux_right_ipin_5.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_right_track_4.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input113_A test_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__281__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mux_right_ipin_3.mux_l2_in_2__A1 sb_1__8_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2__A0 net14 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_10.mux_l2_in_3__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_0__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_11.mux_l4_in_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_83_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_53.mux_l2_in_0_ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_41_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__276__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net239 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_1__A0 sb_1__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net269 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__mux2_4
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input41_A chanx_right_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk sb_1__8_.mem_bottom_track_5.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_1__8_.mem_bottom_track_11.mem_out\[1\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_54_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_11.mux_l3_in_1_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_53.mux_l1_in_1_ net228 net92 sb_1__8_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_11.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_20.mux_l1_in_2__S sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_2.mux_l2_in_1__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_1.mux_l2_in_3_ net341 net232 sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input89_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_43.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_39_prog_clk
+ sb_1__8_.mem_bottom_track_43.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_43.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_23.mux_l1_in_1__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_5.mux_l2_in_1__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_3__252 VGND VGND VPWR VPWR net252 cby_1__8_.mux_right_ipin_1.mux_l2_in_3__252/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_11.mux_l2_in_2_ net232 net230 sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net302 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__284__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_10.ccff_head
+ net239 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_1__8_.mux_bottom_track_9.mux_l1_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ net29 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_17.mux_l2_in_0_ net8 sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_17.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_1.mux_l4_in_0_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sb_1__8_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_left_track_11.mux_l1_in_3_ net228 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_5.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_4.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input106_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input71_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_0__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_3__263 VGND VGND VPWR VPWR net263 cby_1__8_.mux_right_ipin_6.mux_l2_in_3__263/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0__A0 sb_1__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_28.mux_l1_in_3_ net357 net14 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__292__A sb_1__8_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_1.mux_l3_in_1_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_bottom_track_19.mux_l1_in_0__A0 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_80_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__A0 sb_1__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_16_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_2.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ sb_1__8_.mem_bottom_track_11.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input34_A chanx_right_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_4.mux_l2_in_3_ net359 net30 sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_75_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__287__A sb_1__8_.mux_left_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_11.mux_l3_in_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_7_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_53.mux_l1_in_0_ net75 net35 sb_1__8_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_11.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_right_track_2.mux_l2_in_1__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l2_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_1.mux_l2_in_2_ net229 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3__A0 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_43.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk
+ sb_1__8_.mem_bottom_track_41.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_43.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_left_track_5.mux_l2_in_1__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_right_track_28.mux_l3_in_0_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_39_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_11.mux_l2_in_1_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_0.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_1__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk sb_1__8_.mem_bottom_track_17.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_3.mux_l2_in_3__A1 net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_4.mux_l4_in_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_59_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_53.mux_l2_in_1__350 VGND VGND VPWR VPWR net350 sb_1__8_.mux_left_track_53.mux_l2_in_1__350/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_9.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__295__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ net28 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_28.mux_l2_in_1_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk
+ sb_1__8_.mem_bottom_track_49.mem_out\[0\] net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_49.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__274
+ VGND VGND VPWR VPWR net274 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__274/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__8_.mux_left_track_11.mux_l1_in_2_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net87 sb_1__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input64_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_60_prog_clk cby_1__8_.mem_right_ipin_5.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_bottom_track_27.mux_l1_in_0__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_52.mux_l2_in_1__361 VGND VGND VPWR VPWR net361 sb_1__8_.mux_right_track_52.mux_l2_in_1__361/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output220_A net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_4.mux_l3_in_1_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_28.mux_l1_in_2_ net9 net88 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_17.mux_l1_in_0_ net218 net38 sb_1__8_.mem_bottom_track_17.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mux_right_ipin_7.mux_l1_in_2__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_1.mux_l3_in_0_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_19.mux_l1_in_0__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_29.mux_l2_in_0_ net325 sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_29.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_14.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_31.mux_l2_in_0_ net327 sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_31.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_11.ccff_head net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_4.mux_l2_in_2_ net17 net63 sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_0__S sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_9.mux_l2_in_1__340 VGND VGND VPWR VPWR net340 sb_1__8_.mux_bottom_track_9.mux_l2_in_1__340/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_1.mux_l2_in_1__315 VGND VGND VPWR VPWR net315 sb_1__8_.mux_bottom_track_1.mux_l2_in_1__315/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_1.mux_l2_in_1_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net91 sb_1__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_1__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3__A1 net8 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_10_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__298__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 sb_1__8_.mux_bottom_track_25.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_1__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_11.mux_l2_in_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_5.mux_l2_in_3__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input94_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_sb_1__8_.mux_left_track_29.mux_l1_in_1__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_17.mux_l2_in_1__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk cby_1__8_.mem_right_ipin_8.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__286
+ VGND VGND VPWR VPWR net286 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__286/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_1__8_.mem_bottom_track_17.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_17.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_3__258 VGND VGND VPWR VPWR net258 cby_1__8_.mux_right_ipin_15.mux_l2_in_3__258/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_35.mux_l1_in_0__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0__A0 sb_1__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_297_ sb_1__8_.mux_right_track_52.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_28.mux_l2_in_0_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk
+ sb_1__8_.mem_bottom_track_47.ccff_tail net239 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_49.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_2__A0 sb_1__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_left_track_11.mux_l1_in_1_ net69 net81 sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_3__A0 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input1_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_bottom_track_27.mux_l1_in_0__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input57_A chanx_right_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_right_track_4.mux_l3_in_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net283 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_1.mux_l2_in_3__S sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_349_ sb_1__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3_ net370 net62 cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_5.mux_l3_in_0_ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_4__A0 sb_1__8_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_28.mux_l1_in_1_ net70 net82 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input111_A right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_11_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.out sky130_fd_sc_hd__clkbuf_2
XFILLER_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_left_track_7.mux_l2_in_2__A0 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_left_track_45.mux_l1_in_1__A0 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1__A0 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_4.mux_l2_in_1_ net65 net77 sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_3_ net252 sb_1__8_.mux_bottom_track_51.out cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_5.mux_l2_in_1_ net337 net17 sb_1__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net306 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__mux2_4
Xclkbuf_leaf_29_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_1.mux_l2_in_0_ net73 sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_1__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_bottom_track_29.mux_l1_in_0_ net29 net59 sb_1__8_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__298
+ VGND VGND VPWR VPWR net298 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__298/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__8_.mux_left_track_37.mux_l1_in_0__S sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__295
+ VGND VGND VPWR VPWR net295 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__295/LO
+ sky130_fd_sc_hd__conb_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3_ net243 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_43.mux_l1_in_0__A0 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_31.mux_l1_in_0_ net28 net58 sb_1__8_.mem_bottom_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_62_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_6.mux_l1_in_1__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_43.mux_l2_in_0_ net333 sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_43.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input87_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__A1 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__8_.mux_right_ipin_4.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk sb_1__8_.mem_bottom_track_15.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0__A0 sb_1__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__8_.mux_right_ipin_11.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__8_.mux_bottom_track_35.mux_l1_in_0__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_1.mux_l4_in_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_296_ net26 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out net5
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__mux2_1
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mux_right_ipin_2.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_11.mux_l1_in_0_ net58 net43 sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_left_track_7.mux_l1_in_3__A1 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2__A0 sb_1__8_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_3_ net263 sb_1__8_.mux_bottom_track_49.out cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_348_ sb_1__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
X_279_ sb_1__8_.mux_left_track_29.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_53.mux_l1_in_1__A0 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_29.mux_l1_in_3__345 VGND VGND VPWR VPWR net345 sb_1__8_.mux_left_track_29.mux_l1_in_3__345/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_83_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2_ net31 net39 cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_1.mux_l3_in_1_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mux_bottom_track_1.mux_l1_in_0__A0 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_2__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__8_.mux_right_ipin_9.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_28.mux_l1_in_0_ net104 net110 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input104_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_left_track_7.mux_l2_in_2__A1 net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3_ net248 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__245 VGND VGND VPWR VPWR net245 cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__245/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_left_track_13.mux_l1_in_1__S sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_left_track_45.mux_l1_in_1__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_37.mux_l2_in_1__347 VGND VGND VPWR VPWR net347 sb_1__8_.mux_left_track_37.mux_l2_in_1__347/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_4_ sb_1__8_.mux_bottom_track_37.out net65 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_58_prog_clk cby_1__8_.mem_right_ipin_1.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_right_track_4.mux_l2_in_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_2_ net87 sb_1__8_.mux_bottom_track_33.out cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_1__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_bottom_track_51.mux_l1_in_0__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_5.mux_l2_in_0_ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_0.mux_l2_in_3__A1 sb_1__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__S cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_6.mux_l4_in_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_3_ net255 sb_1__8_.mux_bottom_track_49.out
+ cby_1__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_36.mux_l2_in_1__358 VGND VGND VPWR VPWR net358 sb_1__8_.mux_right_track_36.mux_l2_in_1__358/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net237 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_4.mux_l1_in_1_ net107 net104 sb_1__8_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_19_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_bottom_track_5.mux_l1_in_1_ net20 net221 sb_1__8_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_41.mux_l2_in_0__332 VGND VGND VPWR VPWR net332 sb_1__8_.mux_bottom_track_41.mux_l2_in_0__332/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_6.mux_l3_in_1_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3_ net363 net59 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mux_left_track_1.mux_l1_in_0_ net34 net51 sb_1__8_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_4_ sb_1__8_.mux_bottom_track_37.out net65 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net272 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk sb_1__8_.mem_left_track_11.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_23.mux_l1_in_1__322 VGND VGND VPWR VPWR net322 sb_1__8_.mux_bottom_track_23.mux_l1_in_1__322/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net238 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_295_ net25 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net237
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__8_.mux_right_track_36.mux_l1_in_1__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_12.mux_l4_in_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_17_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net238
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_43.mux_l1_in_0_ net219 net36 sb_1__8_.mem_bottom_track_43.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk cby_1__8_.mem_right_ipin_4.ccff_tail
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_2_ net88 cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out
+ net5 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_347_ sb_1__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_278_ net39 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__8_.mux_left_track_53.mux_l1_in_1__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_1.mux_l3_in_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1_ net8 cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_28.mux_l1_in_1__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3__S cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__8_.mux_bottom_track_1.mux_l1_in_0__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput230 net230 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mux_right_track_10.mux_l1_in_0__S sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A chanx_right_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_12.mux_l3_in_1_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__309
+ VGND VGND VPWR VPWR net309 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__309/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2_ net26 net37 cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net236 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__8_.mux_right_ipin_15.mux_l1_in_0__A0 sb_1__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__8_.mux_right_track_4.mux_l2_in_1__S sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net279 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_3_ sb_1__8_.mux_bottom_track_25.out net71 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_28.mux_l1_in_3__357 VGND VGND VPWR VPWR net357 sb_1__8_.mux_right_track_28.mux_l1_in_3__357/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_1_ net67 cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_6.mux_l1_in_1__A0 sb_1__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__8_.mux_left_track_11.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ sb_1__8_.mem_bottom_track_35.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_35.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net239 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_57_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_2_ net88 cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1__A0 sb_1__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net288 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__mux2_4
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__307
+ VGND VGND VPWR VPWR net307 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__307/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 sb_1__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_38_prog_clk sb_1__8_.mem_right_track_52.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_4.mux_l1_in_0_ net101 net110 sb_1__8_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net235 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_1.mux_l1_in_2_ sb_1__8_.mux_bottom_track_15.out net77 cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_13_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__A0 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_right_track_44.mux_l1_in_1__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_5.mux_l1_in_0_ net218 net47 sb_1__8_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_7.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output229_A net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_6.mux_l3_in_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__8_.mux_right_ipin_13.mux_l2_in_1__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__8_.mux_bottom_track_37.mux_l2_in_0__A0 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_3_ sb_1__8_.mux_bottom_track_25.out net71 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
.ends

