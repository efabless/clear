magic
tech sky130A
magscale 1 2
timestamp 1656942844
<< obsli1 >>
rect 1104 2159 18860 14705
<< obsm1 >>
rect 1104 1776 19398 15020
<< metal2 >>
rect 2042 16400 2098 17200
rect 5998 16400 6054 17200
rect 9954 16400 10010 17200
rect 13910 16400 13966 17200
rect 17866 16400 17922 17200
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
<< obsm2 >>
rect 1214 16344 1986 16538
rect 2154 16344 5942 16538
rect 6110 16344 9898 16538
rect 10066 16344 13854 16538
rect 14022 16344 17810 16538
rect 17978 16344 19392 16538
rect 1214 856 19392 16344
rect 1326 734 1986 856
rect 2154 734 2814 856
rect 2982 734 3642 856
rect 3810 734 4470 856
rect 4638 734 5298 856
rect 5466 734 6126 856
rect 6294 734 6954 856
rect 7122 734 7782 856
rect 7950 734 8610 856
rect 8778 734 9438 856
rect 9606 734 10266 856
rect 10434 734 11094 856
rect 11262 734 11922 856
rect 12090 734 12750 856
rect 12918 734 13578 856
rect 13746 734 14406 856
rect 14574 734 15234 856
rect 15402 734 16062 856
rect 16230 734 16890 856
rect 17058 734 17718 856
rect 17886 734 18546 856
rect 18714 734 19392 856
<< metal3 >>
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 0 14832 800 14952
rect 0 14560 800 14680
rect 0 14288 800 14408
rect 0 14016 800 14136
rect 0 13744 800 13864
rect 0 13472 800 13592
rect 0 13200 800 13320
rect 0 12928 800 13048
rect 0 12656 800 12776
rect 0 12384 800 12504
rect 0 12112 800 12232
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 0 11296 800 11416
rect 0 11024 800 11144
rect 0 10752 800 10872
rect 0 10480 800 10600
rect 0 10208 800 10328
rect 0 9936 800 10056
rect 0 9664 800 9784
rect 0 9392 800 9512
rect 0 9120 800 9240
rect 0 8848 800 8968
rect 0 8576 800 8696
rect 0 8304 800 8424
rect 0 8032 800 8152
rect 0 7760 800 7880
rect 0 7488 800 7608
rect 0 7216 800 7336
rect 0 6944 800 7064
rect 0 6672 800 6792
rect 0 6400 800 6520
rect 0 6128 800 6248
rect 0 5856 800 5976
rect 0 5584 800 5704
rect 0 5312 800 5432
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 0 4496 800 4616
rect 0 4224 800 4344
rect 0 3952 800 4072
rect 0 3680 800 3800
rect 0 3408 800 3528
rect 0 3136 800 3256
rect 0 2864 800 2984
rect 0 2592 800 2712
rect 0 2320 800 2440
rect 19200 14424 20000 14544
rect 19200 14152 20000 14272
rect 19200 13880 20000 14000
rect 19200 13608 20000 13728
rect 19200 13336 20000 13456
rect 19200 13064 20000 13184
rect 19200 12792 20000 12912
rect 19200 12520 20000 12640
rect 19200 12248 20000 12368
rect 19200 11976 20000 12096
rect 19200 11704 20000 11824
rect 19200 11432 20000 11552
rect 19200 11160 20000 11280
rect 19200 10888 20000 11008
rect 19200 10616 20000 10736
rect 19200 10344 20000 10464
rect 19200 10072 20000 10192
rect 19200 9800 20000 9920
rect 19200 9528 20000 9648
rect 19200 9256 20000 9376
rect 19200 8984 20000 9104
rect 19200 8712 20000 8832
rect 19200 8440 20000 8560
rect 19200 8168 20000 8288
rect 19200 7896 20000 8016
rect 19200 7624 20000 7744
rect 19200 7352 20000 7472
rect 19200 7080 20000 7200
rect 19200 6808 20000 6928
rect 19200 6536 20000 6656
rect 19200 6264 20000 6384
rect 19200 5992 20000 6112
rect 19200 5720 20000 5840
rect 19200 5448 20000 5568
rect 19200 5176 20000 5296
rect 19200 4904 20000 5024
rect 19200 4632 20000 4752
rect 19200 4360 20000 4480
rect 19200 4088 20000 4208
rect 19200 3816 20000 3936
rect 19200 3544 20000 3664
rect 19200 3272 20000 3392
rect 19200 3000 20000 3120
rect 19200 2728 20000 2848
rect 19200 2456 20000 2576
rect 0 2048 800 2168
rect 0 1776 800 1896
rect 0 1504 800 1624
<< obsm3 >>
rect 880 14624 19200 15469
rect 880 2376 19120 14624
rect 880 1531 19200 2376
<< metal4 >>
rect 3168 2128 3488 14736
rect 5392 2128 5712 14736
rect 7616 2128 7936 14736
rect 9840 2128 10160 14736
rect 12064 2128 12384 14736
rect 14288 2128 14608 14736
rect 16512 2128 16832 14736
<< obsm4 >>
rect 2083 14816 17421 14925
rect 2083 2619 3088 14816
rect 3568 2619 5312 14816
rect 5792 2619 7536 14816
rect 8016 2619 9760 14816
rect 10240 2619 11984 14816
rect 12464 2619 14208 14816
rect 14688 2619 16432 14816
rect 16912 2619 17421 14816
<< labels >>
rlabel metal3 s 0 12656 800 12776 6 REGIN_FEEDTHROUGH
port 1 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 REGOUT_FEEDTHROUGH
port 2 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 SC_IN_BOT
port 3 nsew signal input
rlabel metal2 s 2042 16400 2098 17200 6 SC_IN_TOP
port 4 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 SC_OUT_BOT
port 5 nsew signal output
rlabel metal2 s 5998 16400 6054 17200 6 SC_OUT_TOP
port 6 nsew signal output
rlabel metal4 s 5392 2128 5712 14736 6 VGND
port 7 nsew ground bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VGND
port 7 nsew ground bidirectional
rlabel metal4 s 14288 2128 14608 14736 6 VGND
port 7 nsew ground bidirectional
rlabel metal4 s 3168 2128 3488 14736 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 7616 2128 7936 14736 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 12064 2128 12384 14736 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 16512 2128 16832 14736 6 VPWR
port 8 nsew power bidirectional
rlabel metal2 s 2870 0 2926 800 6 bottom_grid_pin_0_
port 9 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 bottom_grid_pin_10_
port 10 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 bottom_grid_pin_11_
port 11 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 bottom_grid_pin_12_
port 12 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 bottom_grid_pin_13_
port 13 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 bottom_grid_pin_14_
port 14 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 bottom_grid_pin_15_
port 15 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 bottom_grid_pin_1_
port 16 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 bottom_grid_pin_2_
port 17 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 bottom_grid_pin_3_
port 18 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 bottom_grid_pin_4_
port 19 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 bottom_grid_pin_5_
port 20 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 bottom_grid_pin_6_
port 21 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 bottom_grid_pin_7_
port 22 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 bottom_grid_pin_8_
port 23 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_9_
port 24 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 ccff_head
port 25 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 ccff_tail
port 26 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[0]
port 27 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[10]
port 28 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[11]
port 29 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 chanx_left_in[12]
port 30 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[13]
port 31 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[14]
port 32 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 33 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 34 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[17]
port 35 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[18]
port 36 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[19]
port 37 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[1]
port 38 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[2]
port 39 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[3]
port 40 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[4]
port 41 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[5]
port 42 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[6]
port 43 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[7]
port 44 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[8]
port 45 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[9]
port 46 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 chanx_left_out[0]
port 47 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[10]
port 48 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 chanx_left_out[11]
port 49 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 chanx_left_out[12]
port 50 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[13]
port 51 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 chanx_left_out[14]
port 52 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 chanx_left_out[15]
port 53 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 chanx_left_out[16]
port 54 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 chanx_left_out[17]
port 55 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[18]
port 56 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 chanx_left_out[19]
port 57 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[1]
port 58 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 chanx_left_out[2]
port 59 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 chanx_left_out[3]
port 60 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[4]
port 61 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 chanx_left_out[5]
port 62 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 chanx_left_out[6]
port 63 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 64 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 chanx_left_out[8]
port 65 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 chanx_left_out[9]
port 66 nsew signal output
rlabel metal3 s 19200 9256 20000 9376 6 chanx_right_in[0]
port 67 nsew signal input
rlabel metal3 s 19200 11976 20000 12096 6 chanx_right_in[10]
port 68 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 chanx_right_in[11]
port 69 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[12]
port 70 nsew signal input
rlabel metal3 s 19200 12792 20000 12912 6 chanx_right_in[13]
port 71 nsew signal input
rlabel metal3 s 19200 13064 20000 13184 6 chanx_right_in[14]
port 72 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[15]
port 73 nsew signal input
rlabel metal3 s 19200 13608 20000 13728 6 chanx_right_in[16]
port 74 nsew signal input
rlabel metal3 s 19200 13880 20000 14000 6 chanx_right_in[17]
port 75 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[18]
port 76 nsew signal input
rlabel metal3 s 19200 14424 20000 14544 6 chanx_right_in[19]
port 77 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[1]
port 78 nsew signal input
rlabel metal3 s 19200 9800 20000 9920 6 chanx_right_in[2]
port 79 nsew signal input
rlabel metal3 s 19200 10072 20000 10192 6 chanx_right_in[3]
port 80 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 81 nsew signal input
rlabel metal3 s 19200 10616 20000 10736 6 chanx_right_in[5]
port 82 nsew signal input
rlabel metal3 s 19200 10888 20000 11008 6 chanx_right_in[6]
port 83 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[7]
port 84 nsew signal input
rlabel metal3 s 19200 11432 20000 11552 6 chanx_right_in[8]
port 85 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[9]
port 86 nsew signal input
rlabel metal3 s 19200 3816 20000 3936 6 chanx_right_out[0]
port 87 nsew signal output
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[10]
port 88 nsew signal output
rlabel metal3 s 19200 6808 20000 6928 6 chanx_right_out[11]
port 89 nsew signal output
rlabel metal3 s 19200 7080 20000 7200 6 chanx_right_out[12]
port 90 nsew signal output
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[13]
port 91 nsew signal output
rlabel metal3 s 19200 7624 20000 7744 6 chanx_right_out[14]
port 92 nsew signal output
rlabel metal3 s 19200 7896 20000 8016 6 chanx_right_out[15]
port 93 nsew signal output
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[16]
port 94 nsew signal output
rlabel metal3 s 19200 8440 20000 8560 6 chanx_right_out[17]
port 95 nsew signal output
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_out[18]
port 96 nsew signal output
rlabel metal3 s 19200 8984 20000 9104 6 chanx_right_out[19]
port 97 nsew signal output
rlabel metal3 s 19200 4088 20000 4208 6 chanx_right_out[1]
port 98 nsew signal output
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[2]
port 99 nsew signal output
rlabel metal3 s 19200 4632 20000 4752 6 chanx_right_out[3]
port 100 nsew signal output
rlabel metal3 s 19200 4904 20000 5024 6 chanx_right_out[4]
port 101 nsew signal output
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[5]
port 102 nsew signal output
rlabel metal3 s 19200 5448 20000 5568 6 chanx_right_out[6]
port 103 nsew signal output
rlabel metal3 s 19200 5720 20000 5840 6 chanx_right_out[7]
port 104 nsew signal output
rlabel metal3 s 19200 5992 20000 6112 6 chanx_right_out[8]
port 105 nsew signal output
rlabel metal3 s 19200 6264 20000 6384 6 chanx_right_out[9]
port 106 nsew signal output
rlabel metal2 s 9954 16400 10010 17200 6 clk_1_N_out
port 107 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 clk_1_S_out
port 108 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 clk_1_W_in
port 109 nsew signal input
rlabel metal3 s 19200 3544 20000 3664 6 clk_2_E_out
port 110 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 clk_2_W_in
port 111 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 clk_2_W_out
port 112 nsew signal output
rlabel metal3 s 19200 3272 20000 3392 6 clk_3_E_out
port 113 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 clk_3_W_in
port 114 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 clk_3_W_out
port 115 nsew signal output
rlabel metal2 s 13910 16400 13966 17200 6 prog_clk_0_N_in
port 116 nsew signal input
rlabel metal2 s 17866 16400 17922 17200 6 prog_clk_0_W_out
port 117 nsew signal output
rlabel metal3 s 19200 3000 20000 3120 6 prog_clk_1_N_out
port 118 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 prog_clk_1_S_out
port 119 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 prog_clk_1_W_in
port 120 nsew signal input
rlabel metal3 s 19200 2728 20000 2848 6 prog_clk_2_E_out
port 121 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 prog_clk_2_W_in
port 122 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 prog_clk_2_W_out
port 123 nsew signal output
rlabel metal3 s 19200 2456 20000 2576 6 prog_clk_3_E_out
port 124 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 prog_clk_3_W_in
port 125 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 prog_clk_3_W_out
port 126 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 17200
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1136864
string GDS_FILE /home/marwan/clear_signoff_final/openlane/cbx_1__1_/runs/cbx_1__1_/results/signoff/cbx_1__1_.magic.gds
string GDS_START 65030
<< end >>

