magic
tech sky130A
magscale 1 2
timestamp 1625782880
<< obsli1 >>
rect 1104 2159 16008 17425
<< obsm1 >>
rect 198 1708 17006 17944
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1858 19200 1914 20000
rect 2226 19200 2282 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3514 19200 3570 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4802 19200 4858 20000
rect 5170 19200 5226 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6458 19200 6514 20000
rect 6826 19200 6882 20000
rect 7286 19200 7342 20000
rect 7746 19200 7802 20000
rect 8114 19200 8170 20000
rect 8574 19200 8630 20000
rect 8942 19200 8998 20000
rect 9402 19200 9458 20000
rect 9770 19200 9826 20000
rect 10230 19200 10286 20000
rect 10690 19200 10746 20000
rect 11058 19200 11114 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12346 19200 12402 20000
rect 12714 19200 12770 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 14002 19200 14058 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15290 19200 15346 20000
rect 15658 19200 15714 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16946 19200 17002 20000
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< obsm2 >>
rect 314 19144 514 19200
rect 682 19144 974 19200
rect 1142 19144 1342 19200
rect 1510 19144 1802 19200
rect 1970 19144 2170 19200
rect 2338 19144 2630 19200
rect 2798 19144 2998 19200
rect 3166 19144 3458 19200
rect 3626 19144 3918 19200
rect 4086 19144 4286 19200
rect 4454 19144 4746 19200
rect 4914 19144 5114 19200
rect 5282 19144 5574 19200
rect 5742 19144 5942 19200
rect 6110 19144 6402 19200
rect 6570 19144 6770 19200
rect 6938 19144 7230 19200
rect 7398 19144 7690 19200
rect 7858 19144 8058 19200
rect 8226 19144 8518 19200
rect 8686 19144 8886 19200
rect 9054 19144 9346 19200
rect 9514 19144 9714 19200
rect 9882 19144 10174 19200
rect 10342 19144 10634 19200
rect 10802 19144 11002 19200
rect 11170 19144 11462 19200
rect 11630 19144 11830 19200
rect 11998 19144 12290 19200
rect 12458 19144 12658 19200
rect 12826 19144 13118 19200
rect 13286 19144 13486 19200
rect 13654 19144 13946 19200
rect 14114 19144 14406 19200
rect 14574 19144 14774 19200
rect 14942 19144 15234 19200
rect 15402 19144 15602 19200
rect 15770 19144 16062 19200
rect 16230 19144 16430 19200
rect 16598 19144 16890 19200
rect 204 856 17000 19144
rect 314 800 514 856
rect 682 800 974 856
rect 1142 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2262 856
rect 2430 800 2722 856
rect 2890 800 3090 856
rect 3258 800 3550 856
rect 3718 800 4010 856
rect 4178 800 4378 856
rect 4546 800 4838 856
rect 5006 800 5298 856
rect 5466 800 5666 856
rect 5834 800 6126 856
rect 6294 800 6586 856
rect 6754 800 6954 856
rect 7122 800 7414 856
rect 7582 800 7874 856
rect 8042 800 8242 856
rect 8410 800 8702 856
rect 8870 800 9162 856
rect 9330 800 9530 856
rect 9698 800 9990 856
rect 10158 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11278 856
rect 11446 800 11738 856
rect 11906 800 12106 856
rect 12274 800 12566 856
rect 12734 800 13026 856
rect 13194 800 13394 856
rect 13562 800 13854 856
rect 14022 800 14314 856
rect 14482 800 14682 856
rect 14850 800 15142 856
rect 15310 800 15602 856
rect 15770 800 15970 856
rect 16138 800 16430 856
rect 16598 800 16890 856
<< metal3 >>
rect 0 18232 800 18352
rect 16400 17416 17200 17536
rect 0 14968 800 15088
rect 16400 12384 17200 12504
rect 0 11568 800 11688
rect 0 8304 800 8424
rect 16400 7352 17200 7472
rect 0 4904 800 5024
rect 16400 2456 17200 2576
rect 0 1640 800 1760
<< obsm3 >>
rect 880 18152 16400 18325
rect 800 17616 16400 18152
rect 800 17336 16320 17616
rect 800 15168 16400 17336
rect 880 14888 16400 15168
rect 800 12584 16400 14888
rect 800 12304 16320 12584
rect 800 11768 16400 12304
rect 880 11488 16400 11768
rect 800 8504 16400 11488
rect 880 8224 16400 8504
rect 800 7552 16400 8224
rect 800 7272 16320 7552
rect 800 5104 16400 7272
rect 880 4824 16400 5104
rect 800 2656 16400 4824
rect 800 2376 16320 2656
rect 800 1840 16400 2376
rect 880 1667 16400 1840
<< metal4 >>
rect 3443 2128 3763 17456
rect 5941 2128 6261 17456
rect 8440 2128 8760 17456
rect 10939 2128 11259 17456
rect 13437 2128 13757 17456
<< obsm4 >>
rect 3843 2128 5861 17456
rect 6341 2128 8360 17456
rect 8840 2128 10859 17456
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 1 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 ccff_head
port 2 nsew signal input
rlabel metal3 s 16400 12384 17200 12504 6 ccff_tail
port 3 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[0]
port 4 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_in[10]
port 5 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[11]
port 6 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_in[12]
port 7 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_in[13]
port 8 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_in[14]
port 9 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_in[15]
port 10 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[16]
port 11 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_in[17]
port 12 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[18]
port 13 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_in[19]
port 14 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[1]
port 15 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[2]
port 16 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[3]
port 17 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[4]
port 18 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[5]
port 19 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[6]
port 20 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[7]
port 21 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[8]
port 22 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[9]
port 23 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 24 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_out[10]
port 25 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[11]
port 26 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_out[12]
port 27 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_out[13]
port 28 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[14]
port 29 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[15]
port 30 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_out[16]
port 31 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 chany_bottom_out[17]
port 32 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_out[18]
port 33 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_out[19]
port 34 nsew signal output
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 35 nsew signal output
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 36 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_out[3]
port 37 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 38 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[5]
port 39 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[6]
port 40 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[7]
port 41 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_out[8]
port 42 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_out[9]
port 43 nsew signal output
rlabel metal2 s 8942 19200 8998 20000 6 chany_top_in[0]
port 44 nsew signal input
rlabel metal2 s 13174 19200 13230 20000 6 chany_top_in[10]
port 45 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[11]
port 46 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[12]
port 47 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[13]
port 48 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 chany_top_in[14]
port 49 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[15]
port 50 nsew signal input
rlabel metal2 s 15658 19200 15714 20000 6 chany_top_in[16]
port 51 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[17]
port 52 nsew signal input
rlabel metal2 s 16486 19200 16542 20000 6 chany_top_in[18]
port 53 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 54 nsew signal input
rlabel metal2 s 9402 19200 9458 20000 6 chany_top_in[1]
port 55 nsew signal input
rlabel metal2 s 9770 19200 9826 20000 6 chany_top_in[2]
port 56 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[3]
port 57 nsew signal input
rlabel metal2 s 10690 19200 10746 20000 6 chany_top_in[4]
port 58 nsew signal input
rlabel metal2 s 11058 19200 11114 20000 6 chany_top_in[5]
port 59 nsew signal input
rlabel metal2 s 11518 19200 11574 20000 6 chany_top_in[6]
port 60 nsew signal input
rlabel metal2 s 11886 19200 11942 20000 6 chany_top_in[7]
port 61 nsew signal input
rlabel metal2 s 12346 19200 12402 20000 6 chany_top_in[8]
port 62 nsew signal input
rlabel metal2 s 12714 19200 12770 20000 6 chany_top_in[9]
port 63 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 64 nsew signal output
rlabel metal2 s 4802 19200 4858 20000 6 chany_top_out[10]
port 65 nsew signal output
rlabel metal2 s 5170 19200 5226 20000 6 chany_top_out[11]
port 66 nsew signal output
rlabel metal2 s 5630 19200 5686 20000 6 chany_top_out[12]
port 67 nsew signal output
rlabel metal2 s 5998 19200 6054 20000 6 chany_top_out[13]
port 68 nsew signal output
rlabel metal2 s 6458 19200 6514 20000 6 chany_top_out[14]
port 69 nsew signal output
rlabel metal2 s 6826 19200 6882 20000 6 chany_top_out[15]
port 70 nsew signal output
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[16]
port 71 nsew signal output
rlabel metal2 s 7746 19200 7802 20000 6 chany_top_out[17]
port 72 nsew signal output
rlabel metal2 s 8114 19200 8170 20000 6 chany_top_out[18]
port 73 nsew signal output
rlabel metal2 s 8574 19200 8630 20000 6 chany_top_out[19]
port 74 nsew signal output
rlabel metal2 s 1030 19200 1086 20000 6 chany_top_out[1]
port 75 nsew signal output
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 76 nsew signal output
rlabel metal2 s 1858 19200 1914 20000 6 chany_top_out[3]
port 77 nsew signal output
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 78 nsew signal output
rlabel metal2 s 2686 19200 2742 20000 6 chany_top_out[5]
port 79 nsew signal output
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 80 nsew signal output
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[7]
port 81 nsew signal output
rlabel metal2 s 3974 19200 4030 20000 6 chany_top_out[8]
port 82 nsew signal output
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[9]
port 83 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 84 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 85 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 86 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 left_grid_pin_0_
port 87 nsew signal output
rlabel metal3 s 16400 7352 17200 7472 6 prog_clk_0_E_in
port 88 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 right_width_0_height_0__pin_0_
port 89 nsew signal input
rlabel metal3 s 16400 2456 17200 2576 6 right_width_0_height_0__pin_1_lower
port 90 nsew signal output
rlabel metal3 s 16400 17416 17200 17536 6 right_width_0_height_0__pin_1_upper
port 91 nsew signal output
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 92 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 94 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 95 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 96 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17200 20000
string LEFview TRUE
string GDS_FILE /project/openlane/cby_0__1_/runs/cby_0__1_/results/magic/cby_0__1_.gds
string GDS_END 534394
string GDS_START 106416
<< end >>

