* NGSPICE file created from bottom_right_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt bottom_right_tile VGND VPWR ccff_head ccff_head_1 ccff_tail ccff_tail_0 chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23]
+ chanx_left_in[24] chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28]
+ chanx_left_in[29] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23]
+ chanx_left_out[24] chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28]
+ chanx_left_out[29] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[20] chany_top_in[21] chany_top_in[22] chany_top_in[23]
+ chany_top_in[24] chany_top_in[25] chany_top_in[26] chany_top_in[27] chany_top_in[28]
+ chany_top_in[29] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[20] chany_top_out[21] chany_top_out[22] chany_top_out[23]
+ chany_top_out[24] chany_top_out[25] chany_top_out[26] chany_top_out[27] chany_top_out[28]
+ chany_top_out[29] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk
+ prog_reset_top_in reset_top_in test_enable_top_in top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ top_width_0_height_0_subtile_1__pin_inpad_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ top_width_0_height_0_subtile_3__pin_inpad_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_6.mux_l2_in_1_ net188 net25 sb_8__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_20.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_13.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_131_ sb_8__0_.mux_top_track_48.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_8__0_.mem_top_track_4.mem_out\[1\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_114_ net34 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_28.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_49.mux_l2_in_0_ net159 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput86 net86 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput97 net97 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_7.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_51.mux_l2_in_0_ net161 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ cbx_8__0_.cbx_8__0_.ccff_head VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_6.mux_l2_in_0_ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_6.mux_l1_in_1_ net78 net73 sb_8__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_83_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_130_ sb_8__0_.mux_top_track_50.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_ net193 net51 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_8__0_.mem_top_track_4.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_113_ net35 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_8__0_.mem_top_track_26.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_ net45 net31 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput87 net87 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput98 net98 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X net82 VGND VGND VPWR
+ VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_8__0_.mem_top_track_40.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_33.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_18.mux_l2_in_0_ sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_20.mux_l2_in_0_ net171 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_20.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_49.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net48 sb_8__0_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_51.mux_l1_in_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
+ net49 sb_8__0_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_6.mux_l1_in_0_ net70 net75 sb_8__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_18.mux_l1_in_1_ net169 net31 sb_8__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_ net25 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_8__0_.mem_top_track_2.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_112_ net36 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_5.mux_l2_in_0_ net160 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_ sb_8__0_.mux_left_track_31.out net8
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.out sky130_fd_sc_hd__clkbuf_2
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput88 net88 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput99 net99 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk sb_8__0_.mem_top_track_38.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_31.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.out sky130_fd_sc_hd__clkbuf_1
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_46.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_18.mux_l1_in_0_ net80 net70 sb_8__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_20.mux_l1_in_0_ net32 net71 sb_8__0_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_top_track_32.mux_l2_in_0_ net177 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_111_ sb_8__0_.mux_left_track_29.out VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_8 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_ sb_8__0_.mux_left_track_19.out net15
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput89 net89 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_5.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net44 sb_8__0_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_6.mux_l2_in_1__188 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.mux_l2_in_1__188/HI
+ net188 sky130_fd_sc_hd__conb_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net63 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xsb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_8__0_.mem_top_track_14.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_4.mux_l2_in_1__181 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.mux_l2_in_1__181/HI
+ net181 sky130_fd_sc_hd__conb_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_44.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_20.mux_l2_in_0__171 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.mux_l2_in_0__171/HI
+ net171 sky130_fd_sc_hd__conb_1
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_110_ sb_8__0_.mux_left_track_31.out VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_8__0_.mem_left_track_51.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_32.mux_l1_in_0_ net9 net79 sb_8__0_.mem_top_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_ sb_8__0_.mux_left_track_7.out net21
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_19.mux_l2_in_0_ net151 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_44.mux_l2_in_0_ sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_4_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_36.mux_l2_in_0__179 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.mux_l2_in_0__179/HI
+ net179 sky130_fd_sc_hd__conb_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_44.mux_l1_in_1_ net184 net16 sb_8__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_8__0_.mem_top_track_12.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_18.mux_l1_in_1__169 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.mux_l1_in_1__169/HI
+ net169 sky130_fd_sc_hd__conb_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193/HI
+ net193 sky130_fd_sc_hd__conb_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_48.mux_l1_in_1__186 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.mux_l1_in_1__186/HI
+ net186 sky130_fd_sc_hd__conb_1
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net66 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.out sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_8__0_.mem_left_track_49.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_ sb_8__0_.mux_left_track_1.out net24
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_19.mux_l1_in_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
+ net61 sb_8__0_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_44.mux_l1_in_0_ net77 net71 sb_8__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_left_track_33.mux_l2_in_0_ net155 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_33.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_2.mux_l3_in_0_ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_099_ net50 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.out sky130_fd_sc_hd__clkbuf_1
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_2.mux_l2_in_1_ net170 net3 sb_8__0_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_8__0_.mem_top_track_32.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_51.mux_l2_in_0__161 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.mux_l2_in_0__161/HI
+ net161 sky130_fd_sc_hd__conb_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_17.mux_l2_in_0__198 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.mux_l2_in_0__198/HI
+ net198 sky130_fd_sc_hd__conb_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_9.mux_l2_in_0__163 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.mux_l2_in_0__163/HI
+ net163 sky130_fd_sc_hd__conb_1
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_33.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net39 sb_8__0_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_45.mux_l2_in_0_ net157 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_098_ net51 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_left_track_35.mux_l2_in_0__156 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.mux_l2_in_0__156/HI
+ net156 sky130_fd_sc_hd__conb_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_2.mux_l2_in_0_ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_8__0_.mem_top_track_30.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_2.mux_l1_in_1_ net79 net74 sb_8__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_13_0_prog_clk cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ net68 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk sb_8__0_.mem_top_track_38.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_38.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_097_ net52 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_14.mux_l2_in_0_ sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_149_ sb_8__0_.mux_top_track_12.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_45.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net46 sb_8__0_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_2.mux_l1_in_0_ net71 net76 sb_8__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_14.mux_l1_in_1_ net167 net29 sb_8__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_53_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_8__0_.mem_top_track_36.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_38.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_1.mux_l2_in_0_ sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_8__0_.mem_top_track_50.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.out sky130_fd_sc_hd__clkbuf_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_1.mux_l1_in_1_ net194 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_096_ net53 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_148_ sb_8__0_.mux_top_track_14.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_14.mux_l1_in_0_ net78 net76 sb_8__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_26.mux_l2_in_0_ net174 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_26.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191/HI
+ net191 sky130_fd_sc_hd__conb_1
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_49.mux_l2_in_0__159 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.mux_l2_in_0__159/HI
+ net159 sky130_fd_sc_hd__conb_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_11.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_89_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_8__0_.mem_top_track_48.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_1.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net54 sb_8__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.out sky130_fd_sc_hd__clkbuf_1
X_147_ sb_8__0_.mux_top_track_16.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_7.mux_l1_in_1__162 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.mux_l1_in_1__162/HI
+ net162 sky130_fd_sc_hd__conb_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_5.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_49.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_34.mux_l2_in_0__178 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.mux_l2_in_0__178/HI
+ net178 sky130_fd_sc_hd__conb_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_2.mux_l2_in_1__170 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.mux_l2_in_1__170/HI
+ net170 sky130_fd_sc_hd__conb_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_16.mux_l1_in_1__168 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.mux_l1_in_1__168/HI
+ net168 sky130_fd_sc_hd__conb_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_26.mux_l1_in_0_ net6 net74 sb_8__0_.mem_top_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_46.mux_l1_in_1__185 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.mux_l1_in_1__185/HI
+ net185 sky130_fd_sc_hd__conb_1
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_11.ccff_head
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_38.mux_l2_in_0_ net180 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_38.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_15.mux_l2_in_0_ net197 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_15.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_40.mux_l2_in_0_ net182 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_8__0_.mem_top_track_0.mem_out\[1\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_163_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_24.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_146_ sb_8__0_.mux_top_track_18.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_17.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_29.mux_l2_in_0__152 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.mux_l2_in_0__152/HI
+ net152 sky130_fd_sc_hd__conb_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_129_ net20 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_47.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_8__0_.mem_left_track_3.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_50.mux_l1_in_1__187 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.mux_l1_in_1__187/HI
+ net187 sky130_fd_sc_hd__conb_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.out sky130_fd_sc_hd__clkbuf_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_top_track_0.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_162_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_8__0_.mem_top_track_22.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_38.mux_l1_in_0_ net12 net76 sb_8__0_.mem_top_track_38.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk net199 VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_15.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net59 sb_8__0_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_145_ sb_8__0_.mux_top_track_20.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_40.mux_l1_in_0_ net13 net69 sb_8__0_.mem_top_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_15.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_128_ net21 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_8__0_.mem_top_track_6.mem_out\[1\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput70 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net70 sky130_fd_sc_hd__buf_2
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_15.mux_l2_in_0__197 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.mux_l2_in_0__197/HI
+ net197 sky130_fd_sc_hd__conb_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk net2
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_161_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_33.mux_l2_in_0__155 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.mux_l2_in_0__155/HI
+ net155 sky130_fd_sc_hd__conb_1
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 ccff_head_1 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_144_ sb_8__0_.mux_top_track_22.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_127_ net22 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_8__0_.mem_top_track_6.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput60 chany_top_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
Xinput71 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net71 sky130_fd_sc_hd__buf_2
XFILLER_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_10.mux_l3_in_0_ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_8__0_.mem_top_track_10.mem_out\[1\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mux_top_track_8.mux_l3_in_0_ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_8__0_.mem_top_track_42.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_42.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_10.mux_l2_in_1_ net165 net27 sb_8__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_35.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_160_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_8.mux_l2_in_1_ net189 net26 sb_8__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_143_ sb_8__0_.mux_top_track_24.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_126_ net23 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_8__0_.mem_top_track_4.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput72 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net72 sky130_fd_sc_hd__buf_2
Xinput50 chany_top_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput61 chany_top_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_109_ sb_8__0_.mux_left_track_33.out VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_8__0_.mem_top_track_10.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_8__0_.mem_top_track_40.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_42.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net81 net67 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_10.mux_l2_in_0_ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_33.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_ net190 sb_8__0_.mux_left_track_49.out
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_8.mux_l2_in_0_ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_10.mux_l1_in_1_ net80 net77 sb_8__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_142_ sb_8__0_.mux_top_track_26.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_48.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_ net41 net5 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_8.mux_l1_in_1_ net79 net74 sb_8__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_125_ sb_8__0_.mux_left_track_1.out VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput40 chany_top_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput73 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net73 sky130_fd_sc_hd__buf_2
Xinput62 chany_top_in[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
Xinput51 chany_top_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_108_ sb_8__0_.mux_left_track_35.out VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_8__0_.mem_top_track_10.ccff_head
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_28.mux_l2_in_0__175 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.mux_l2_in_0__175/HI
+ net175 sky130_fd_sc_hd__conb_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_47.mux_l2_in_0__158 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.mux_l2_in_0__158/HI
+ net158 sky130_fd_sc_hd__conb_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net64 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_16.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail net67
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_10.mux_l1_in_0_ net72 net69 sb_8__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_4_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_46.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_141_ sb_8__0_.mux_top_track_28.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_22.mux_l2_in_0_ net172 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_22.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_ net35 net11 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_21 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput150 net150 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
Xsb_8__0_.mux_top_track_8.mux_l1_in_0_ net71 net76 sb_8__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ sb_8__0_.mux_left_track_3.out VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput52 chany_top_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chany_top_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput63 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net74 sky130_fd_sc_hd__buf_2
Xsb_8__0_.mux_top_track_32.mux_l2_in_0__177 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.mux_l2_in_0__177/HI
+ net177 sky130_fd_sc_hd__conb_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_107_ net41 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_14.mux_l1_in_1__167 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.mux_l1_in_1__167/HI
+ net167 sky130_fd_sc_hd__conb_1
XFILLER_93_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_7.mux_l2_in_0_ sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_left_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_44.mux_l1_in_1__184 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.mux_l1_in_1__184/HI
+ net184 sky130_fd_sc_hd__conb_1
XFILLER_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_7.mux_l1_in_1_ net162 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_8__0_.mem_top_track_14.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.out sky130_fd_sc_hd__clkbuf_1
XFILLER_41_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_140_ sb_8__0_.mux_top_track_30.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_ sb_8__0_.mux_left_track_13.out net18
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_7_0_prog_clk cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ net68 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.out sky130_fd_sc_hd__clkbuf_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput140 net140 VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_123_ sb_8__0_.mux_left_track_5.out VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 chany_top_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 chany_top_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xinput64 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR VPWR
+ net75 sky130_fd_sc_hd__buf_2
XFILLER_88_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_22.mux_l1_in_0_ net4 net72 sb_8__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_34.mux_l2_in_0_ net178 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ net42 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_11.mux_l2_in_0_ net195 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_89_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_5.mux_l2_in_0__160 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.mux_l2_in_0__160/HI
+ net160 sky130_fd_sc_hd__conb_1
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.out sky130_fd_sc_hd__clkbuf_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_7.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net55 sb_8__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_ sb_8__0_.mux_left_track_7.out net21
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_23 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_top_out[25] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_8__0_.mux_left_track_7.out VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput43 chany_top_in[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput54 chany_top_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xinput76 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR VPWR
+ net76 sky130_fd_sc_hd__buf_2
Xinput65 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_105_ net43 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_13.mux_l2_in_0__196 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.mux_l2_in_0__196/HI
+ net196 sky130_fd_sc_hd__conb_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_8__0_.mem_top_track_34.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_34.mux_l1_in_0_ net10 net80 sb_8__0_.mem_top_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_11.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net57 sb_8__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_top_track_46.mux_l2_in_0_ sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_46.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_31.mux_l2_in_0__154 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.mux_l2_in_0__154/HI
+ net154 sky130_fd_sc_hd__conb_1
XFILLER_1_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_46.mux_l1_in_1_ net185 net17 sb_8__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ sb_8__0_.mux_left_track_1.out net24
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_24 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_top_out[26] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_121_ sb_8__0_.mux_left_track_9.out VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 chany_top_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput44 chany_top_in[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput33 chany_top_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput66 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net77 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_104_ net45 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.out sky130_fd_sc_hd__clkbuf_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_32.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_10.mux_l2_in_1__165 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.mux_l2_in_1__165/HI
+ net165 sky130_fd_sc_hd__conb_1
Xsb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_46.mux_l1_in_0_ net78 net72 sb_8__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_35.mux_l2_in_0_ net156 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_35.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_14 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_25 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput110 net110 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chany_top_out[27] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ sb_8__0_.mux_left_track_11.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_top_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 chany_top_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 chany_top_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
Xinput78 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net78 sky130_fd_sc_hd__buf_2
Xinput67 isol_n VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.mux_l3_in_0_ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_103_ sb_8__0_.mux_left_track_45.out VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.mux_l2_in_1_ net181 net14 sb_8__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.out sky130_fd_sc_hd__clkbuf_1
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_26 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput100 net100 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chany_top_out[28] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_top_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_top_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput68 prog_reset_top_in VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_16
Xinput57 chany_top_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput79 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_1.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_45.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_102_ sb_8__0_.mux_left_track_47.out VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_35.mux_l1_in_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
+ net40 sb_8__0_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_47.mux_l2_in_0_ net158 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_26.mux_l2_in_0__174 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.mux_l2_in_0__174/HI
+ net174 sky130_fd_sc_hd__conb_1
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.mux_l2_in_0_ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_45.mux_l2_in_0__157 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.mux_l2_in_0__157/HI
+ net157 sky130_fd_sc_hd__conb_1
XFILLER_74_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_4.mux_l1_in_1_ net80 net77 sb_8__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_81_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_20.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_ net191 sb_8__0_.mux_left_track_51.out
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_27 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_13.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chany_top_out[29] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_top_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput69 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net69 sky130_fd_sc_hd__buf_2
Xinput47 chany_top_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 chany_top_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_30.mux_l2_in_0__176 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.mux_l2_in_0__176/HI
+ net176 sky130_fd_sc_hd__conb_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_8__0_.mem_left_track_1.ccff_head
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_35.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_ net42 net4 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_101_ sb_8__0_.mux_left_track_49.out VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_0.mux_l2_in_1__164 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.mux_l2_in_1__164/HI
+ net164 sky130_fd_sc_hd__conb_1
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_12.mux_l1_in_1__166 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.mux_l1_in_1__166/HI
+ net166 sky130_fd_sc_hd__conb_1
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_16.mux_l2_in_0_ sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_8__0_.mem_left_track_7.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_47.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net47 sb_8__0_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.mux_l1_in_0_ net72 net69 sb_8__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_16.mux_l1_in_1_ net168 net30 sb_8__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_18.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xwire1 prog_clk VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_ net27 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_11.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_12
Xoutput102 net102 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_3.mux_l2_in_0_ net153 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 chany_top_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput59 chany_top_in[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput48 chany_top_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_38.mux_l2_in_0__180 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.mux_l2_in_0__180/HI
+ net180 sky130_fd_sc_hd__conb_1
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_8__0_.mem_top_track_2.mem_out\[1\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_ net36 net10 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.out sky130_fd_sc_hd__clkbuf_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_100_ sb_8__0_.mux_left_track_51.out VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_26.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_19.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_8__0_.mem_left_track_5.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_16.mux_l1_in_0_ net79 net69 sb_8__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_28.mux_l2_in_0_ net175 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_30.mux_l2_in_0_ net176 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chany_top_out[20] sky130_fd_sc_hd__buf_12
Xoutput103 net103 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 chany_top_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput49 chany_top_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_8__0_.mem_top_track_2.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_ sb_8__0_.mux_left_track_15.out net17
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_24.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_11.mux_l2_in_0__195 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.mux_l2_in_0__195/HI
+ net195 sky130_fd_sc_hd__conb_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_159_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_3.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net33 sb_8__0_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_8__0_.mem_left_track_17.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_8__0_.mem_top_track_8.mem_out\[1\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.out sky130_fd_sc_hd__clkbuf_1
XFILLER_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_31.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192/HI
+ net192 sky130_fd_sc_hd__conb_1
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_42.mux_l2_in_0__183 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.mux_l2_in_0__183/HI
+ net183 sky130_fd_sc_hd__conb_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_1
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_19 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput115 net115 VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_12
Xoutput104 net104 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chany_top_out[21] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput39 chany_top_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_28.mux_l1_in_0_ net7 net77 sb_8__0_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_8__0_.mem_top_track_0.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_30.mux_l1_in_0_ net8 net78 sb_8__0_.mem_top_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_ sb_8__0_.mux_left_track_9.out net20
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_17.mux_l2_in_0_ net198 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_17.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_42.mux_l2_in_0_ net183 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_158_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_8__0_.mem_top_track_8.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_29.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_8__0_.mem_top_track_44.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput138 net138 VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_top_out[22] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
XFILLER_95_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_ sb_8__0_.mux_left_track_3.out net23
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_157_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_17.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net60 sb_8__0_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_8__0_.mem_top_track_6.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_42.mux_l1_in_0_ net15 net70 sb_8__0_.mem_top_track_42.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_79_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_29.mux_l2_in_0_ net152 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_29.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_4_0_prog_clk net1 net68 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_31.mux_l2_in_0_ net154 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_31.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_12.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_0.mux_l3_in_0_ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_8__0_.mem_top_track_42.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput106 net106 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_top_out[23] sky130_fd_sc_hd__buf_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_0.mux_l2_in_1_ net164 net24 sb_8__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_156_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_24.mux_l2_in_0__173 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.mux_l2_in_0__173/HI
+ net173 sky130_fd_sc_hd__conb_1
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_139_ sb_8__0_.mux_top_track_32.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_88_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_5_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_10.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_29.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net37 sb_8__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_31.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net38 sb_8__0_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput107 net107 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_top_out[24] sky130_fd_sc_hd__buf_12
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net65 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_77_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_0.mux_l2_in_0_ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_8__0_.mem_top_track_18.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_155_ sb_8__0_.mux_top_track_0.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_8_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\] net68 VGND VGND VPWR VPWR net82
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_3.mux_l2_in_0__153 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.mux_l2_in_0__153/HI
+ net153 sky130_fd_sc_hd__conb_1
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_0.mux_l1_in_1_ net78 net73 sb_8__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_138_ sb_8__0_.mux_top_track_34.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput119 net119 VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_12
Xoutput108 net108 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput90 net90 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
XFILLER_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_16.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_12.mux_l2_in_0_ sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_ net192 net50 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_154_ sb_8__0_.mux_top_track_2.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_0.mux_l1_in_0_ net70 net75 sb_8__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_8__0_.mem_top_track_30.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_12.mux_l1_in_1_ net166 net28 sb_8__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_137_ sb_8__0_.mux_top_track_36.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_ net43 net32 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190/HI
+ net190 sky130_fd_sc_hd__conb_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net109 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput91 net91 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
XFILLER_95_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_1.mux_l1_in_1__194 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.mux_l1_in_1__194/HI
+ net194 sky130_fd_sc_hd__conb_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ sb_8__0_.mux_top_track_4.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_77_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_8__0_.mem_top_track_28.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_12.mux_l1_in_0_ net77 net75 sb_8__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_136_ sb_8__0_.mux_top_track_38.out VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_24.mux_l2_in_0_ net173 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_24.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_ sb_8__0_.mux_left_track_29.out net9
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk
+ cbx_8__0_.cbx_8__0_.ccff_head net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_119_ sb_8__0_.mux_left_track_13.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_8__0_.mem_top_track_36.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_40.mux_l2_in_0__182 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.mux_l2_in_0__182/HI
+ net182 sky130_fd_sc_hd__conb_1
XFILLER_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_29.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput92 net92 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput81 net81 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XFILLER_95_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_9.mux_l2_in_0_ net163 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.out sky130_fd_sc_hd__clkbuf_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_152_ sb_8__0_.mux_top_track_6.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail net68 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_26_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_135_ sb_8__0_.mux_top_track_40.out VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_ sb_8__0_.mux_left_track_17.out net16
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_118_ sb_8__0_.mux_left_track_15.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.out sky130_fd_sc_hd__clkbuf_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_24.mux_l1_in_0_ net5 net73 sb_8__0_.mem_top_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_8__0_.mem_top_track_34.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_36.mux_l2_in_0_ net179 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_36.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_13.mux_l2_in_0_ net196 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_19.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput93 net93 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_19.mux_l2_in_0__151 VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.mux_l2_in_0__151/HI
+ net151 sky130_fd_sc_hd__conb_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_151_ sb_8__0_.mux_top_track_8.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_9.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net56 sb_8__0_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_134_ sb_8__0_.mux_top_track_42.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_ sb_8__0_.mux_left_track_11.out net19
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.out sky130_fd_sc_hd__clkbuf_1
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ sb_8__0_.mux_left_track_17.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput83 net83 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput94 net94 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail net67
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xsb_8__0_.mux_top_track_36.mux_l1_in_0_ net11 net75 sb_8__0_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_8.mux_l2_in_1__189 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.mux_l2_in_1__189/HI
+ net189 sky130_fd_sc_hd__conb_1
Xsb_8__0_.mux_left_track_13.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net58 sb_8__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_48.mux_l2_in_0_ sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_48.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_150_ sb_8__0_.mux_top_track_10.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_50.mux_l2_in_0_ sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_left_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_22.mux_l2_in_0__172 VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.mux_l2_in_0__172/HI
+ net172 sky130_fd_sc_hd__conb_1
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_13_0_prog_clk cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ net68 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfrtp_4
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_133_ sb_8__0_.mux_top_track_44.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_48.mux_l1_in_1_ net186 net18 sb_8__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_ sb_8__0_.mux_left_track_5.out net22
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_50.mux_l1_in_1_ net187 net19 sb_8__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_47.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_8__0_.mem_left_track_3.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_116_ sb_8__0_.mux_left_track_19.out VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput84 net84 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput95 net95 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
XFILLER_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.out sky130_fd_sc_hd__clkbuf_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_8__0_.mem_top_track_22.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail net67
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_15.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_132_ sb_8__0_.mux_top_track_46.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_48.mux_l1_in_0_ net79 net73 sb_8__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_50.mux_l1_in_0_ net80 net74 sb_8__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_8__0_.mem_left_track_1.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_8__0_.mem_left_track_45.ccff_tail
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ net62 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_6.mux_l3_in_0_ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput85 net85 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput96 net96 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
XFILLER_48_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_8__0_.mem_left_track_9.mem_out\[0\]
+ net68 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

